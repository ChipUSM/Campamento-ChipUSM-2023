magic
tech sky130A
timestamp 1702349019
<< error_p >>
rect -166 181 166 183
rect -166 -181 -151 181
rect -133 148 133 150
rect -133 -148 -118 148
rect 118 -148 133 148
rect -133 -150 133 -148
rect 151 -181 166 181
rect -166 -183 166 -181
<< nwell >>
rect -151 -181 151 181
<< mvpmos >>
rect -104 -150 -54 150
rect -25 -150 25 150
rect 54 -150 104 150
<< mvpdiff >>
rect -133 144 -104 150
rect -133 -144 -127 144
rect -110 -144 -104 144
rect -133 -150 -104 -144
rect -54 144 -25 150
rect -54 -144 -48 144
rect -31 -144 -25 144
rect -54 -150 -25 -144
rect 25 144 54 150
rect 25 -144 31 144
rect 48 -144 54 144
rect 25 -150 54 -144
rect 104 144 133 150
rect 104 -144 110 144
rect 127 -144 133 144
rect 104 -150 133 -144
<< mvpdiffc >>
rect -127 -144 -110 144
rect -48 -144 -31 144
rect 31 -144 48 144
rect 110 -144 127 144
<< poly >>
rect -104 150 -54 163
rect -25 150 25 163
rect 54 150 104 163
rect -104 -163 -54 -150
rect -25 -163 25 -150
rect 54 -163 104 -150
<< locali >>
rect -127 144 -110 152
rect -127 -152 -110 -144
rect -48 144 -31 152
rect -48 -152 -31 -144
rect 31 144 48 152
rect 31 -152 48 -144
rect 110 144 127 152
rect 110 -152 127 -144
<< viali >>
rect -127 -144 -110 144
rect -48 -144 -31 144
rect 31 -144 48 144
rect 110 -144 127 144
<< metal1 >>
rect -130 144 -107 150
rect -130 -144 -127 144
rect -110 -144 -107 144
rect -130 -150 -107 -144
rect -51 144 -28 150
rect -51 -144 -48 144
rect -31 -144 -28 144
rect -51 -150 -28 -144
rect 28 144 51 150
rect 28 -144 31 144
rect 48 -144 51 144
rect 28 -150 51 -144
rect 107 144 130 150
rect 107 -144 110 144
rect 127 -144 130 144
rect 107 -150 130 -144
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 3 l 0.5 m 1 nf 3 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
