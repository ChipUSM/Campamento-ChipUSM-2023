magic
tech sky130A
magscale 1 2
timestamp 1702647744
<< error_p >>
rect 8222 5114 8238 5130
rect 9362 5114 9378 5130
rect 8206 5098 8222 5114
rect 9378 5098 9394 5114
rect 8221 4166 9376 4172
rect 346 3800 1236 3836
rect 346 3000 382 3800
rect 1200 3000 1236 3800
rect 346 2964 1236 3000
rect 1964 3800 2854 3836
rect 1964 3000 2000 3800
rect 2818 3000 2854 3800
rect 8221 3788 8227 4166
rect 9370 3170 9376 4166
rect 9118 3164 9376 3170
rect 1964 2964 2854 3000
rect 8206 2959 8222 2975
rect 9378 2959 9394 2975
rect 8222 2943 8238 2959
rect 9362 2943 9378 2959
rect 800 1400 816 1416
rect 1584 1400 1600 1416
rect 2400 1400 2416 1416
rect 3184 1400 3200 1416
rect 784 1384 808 1400
rect 1600 1384 1616 1400
rect 2384 1384 2400 1400
rect 3200 1384 3216 1400
rect 800 616 808 1384
rect 784 608 808 616
rect 1600 608 1616 616
rect 784 600 1616 608
rect 2384 608 2400 616
rect 3200 608 3216 616
rect 2384 600 3216 608
rect 800 584 816 600
rect 1584 584 1600 600
rect 2400 584 2416 600
rect 3184 584 3200 600
rect 800 -1400 816 -1384
rect 1584 -1400 1600 -1384
rect 2400 -1400 2416 -1384
rect 3184 -1400 3200 -1384
rect 784 -1408 1616 -1400
rect 784 -1416 808 -1408
rect 1600 -1416 1616 -1408
rect 2384 -1408 3216 -1400
rect 2384 -1416 2400 -1408
rect 3200 -1416 3216 -1408
rect 800 -2184 808 -1416
rect 784 -2200 808 -2184
rect 1600 -2200 1616 -2184
rect 2384 -2200 2400 -2184
rect 3200 -2200 3216 -2184
rect 800 -2216 816 -2200
rect 1584 -2216 1600 -2200
rect 2400 -2216 2416 -2200
rect 3184 -2216 3200 -2200
rect 400 -3400 424 -3376
rect 1176 -3400 1200 -3376
rect 2000 -3400 2024 -3376
rect 2776 -3400 2800 -3376
rect 376 -3424 400 -3400
rect 1200 -3424 1224 -3400
rect 1976 -3424 2000 -3400
rect 2800 -3424 2824 -3400
rect 376 -4200 400 -4176
rect 1200 -4200 1224 -4176
rect 1976 -4200 2000 -4176
rect 2800 -4200 2824 -4176
rect 400 -4224 424 -4200
rect 1176 -4224 1200 -4200
rect 2000 -4224 2024 -4200
rect 2776 -4224 2800 -4200
<< nwell >>
rect 7059 2430 10423 5565
rect 0 0 4000 2200
<< nmos >>
rect 1800 -2400 2200 -1400
<< pmos >>
rect 1800 600 2200 1600
<< ndiff >>
rect 1600 -2200 1800 -1400
rect 800 -2400 1800 -2200
rect 2200 -2200 2400 -1400
rect 3200 -2200 3400 -1400
rect 2200 -2400 3400 -2200
<< pdiff >>
rect 800 1400 1800 1600
rect 1600 600 1800 1400
rect 2200 1400 3400 1600
rect 2200 600 2400 1400
rect 3200 600 3400 1400
<< ndiffc >>
rect 800 -2200 1600 -1400
rect 2400 -2200 3200 -1400
<< pdiffc >>
rect 800 600 1600 1400
rect 2400 600 3200 1400
<< nsubdiff >>
rect 7672 5114 9919 5169
rect 7672 2959 8222 5114
rect 9378 2959 9919 5114
rect 7672 2904 9919 2959
<< psubdiffcont >>
rect 400 -4200 1200 -3400
rect 2000 -4200 2800 -3400
<< nsubdiffcont >>
rect 382 3000 1200 3800
rect 2000 3000 2818 3800
rect 8222 2959 9378 5114
<< poly >>
rect 1800 1600 2200 2000
rect 1800 -200 2200 600
rect 1400 -1000 2200 -200
rect 1800 -1400 2200 -1000
rect 1800 -2800 2200 -2400
<< viali >>
rect 8221 3164 8222 4172
rect 8222 3164 9376 4172
<< metal1 >>
rect 400 3794 3400 3800
rect 400 3164 8221 3794
rect 400 3000 9124 3164
rect 800 600 1600 3000
rect 3299 2965 9124 3000
rect 2400 -200 3200 1400
rect 2400 -1000 4000 -200
rect 800 -3400 1600 -1400
rect 2400 -2200 3200 -1000
rect 400 -4200 3600 -3400
<< labels >>
rlabel metal1 3200 -800 3400 -600 1 out
port 1 n
rlabel poly 1600 -800 1800 -600 1 in
port 2 n
rlabel metal1 1200 -3800 1400 -3600 1 gnd
port 3 n
rlabel metal1 1200 3400 1400 3600 1 vdd
port 4 n
<< end >>
