magic
tech sky130A
magscale 1 2
timestamp 1702349019
<< error_p >>
rect -253 112 253 116
rect -253 -112 -223 112
rect -187 46 187 50
rect -187 -46 -157 46
rect 157 -46 187 46
rect -187 -50 187 -46
rect 223 -112 253 112
rect -253 -116 253 -112
<< nwell >>
rect -223 -112 223 112
<< mvpmos >>
rect -129 -50 -29 50
rect 29 -50 129 50
<< mvpdiff >>
rect -187 38 -129 50
rect -187 -38 -175 38
rect -141 -38 -129 38
rect -187 -50 -129 -38
rect -29 38 29 50
rect -29 -38 -17 38
rect 17 -38 29 38
rect -29 -50 29 -38
rect 129 38 187 50
rect 129 -38 141 38
rect 175 -38 187 38
rect 129 -50 187 -38
<< mvpdiffc >>
rect -175 -38 -141 38
rect -17 -38 17 38
rect 141 -38 175 38
<< poly >>
rect -129 50 -29 76
rect 29 50 129 76
rect -129 -76 -29 -50
rect 29 -76 129 -50
<< locali >>
rect -175 38 -141 54
rect -175 -54 -141 -38
rect -17 38 17 54
rect -17 -54 17 -38
rect 141 38 175 54
rect 141 -54 175 -38
<< viali >>
rect -175 -38 -141 38
rect -17 -38 17 38
rect 141 -38 175 38
<< metal1 >>
rect -181 38 -135 50
rect -181 -38 -175 38
rect -141 -38 -135 38
rect -181 -50 -135 -38
rect -23 38 23 50
rect -23 -38 -17 38
rect 17 -38 23 38
rect -23 -50 23 -38
rect 135 38 181 50
rect 135 -38 141 38
rect 175 -38 181 38
rect 135 -50 181 -38
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 0.5 l 0.5 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
