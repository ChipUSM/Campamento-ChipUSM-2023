magic
tech sky130A
magscale 1 2
timestamp 1702583177
<< dnwell >>
rect -1650 2992 -856 3602
rect -1650 42 -856 652
rect -1650 -2912 -856 -2302
<< nwell >>
rect -1720 5322 -632 5538
rect -1720 5206 -768 5322
rect -1720 3714 -1552 5206
rect -1274 4502 -768 5206
rect -1720 3546 -822 3714
rect -1720 3144 -1508 3546
rect -990 3144 -822 3546
rect -1720 2980 -822 3144
rect -1722 2976 -822 2980
rect -1722 2588 -824 2976
rect -1722 2586 -632 2588
rect -1720 2372 -632 2586
rect 1408 2562 1914 2616
rect 2308 2562 2814 2616
rect 3258 2590 3718 2658
rect -1720 2256 -768 2372
rect 1408 2344 2050 2562
rect 2308 2344 2950 2562
rect 3204 2362 3718 2590
rect 3206 2346 3718 2362
rect 1408 2284 1914 2344
rect 2308 2284 2814 2344
rect 3370 2316 3718 2346
rect -1720 764 -1552 2256
rect -1274 1552 -768 2256
rect 420 2046 926 2100
rect 420 1828 1062 2046
rect 420 1768 926 1828
rect 1408 1660 1914 1714
rect 1408 1442 2050 1660
rect 2304 1504 2810 1558
rect 3258 1532 3718 1600
rect 1408 1382 1914 1442
rect 2304 1282 2946 1504
rect 3204 1304 3718 1532
rect 3206 1288 3718 1304
rect 2304 1226 2822 1282
rect 3370 1258 3718 1288
rect -1720 596 -822 764
rect -1720 194 -1508 596
rect -990 194 -822 596
rect 420 698 926 752
rect 1372 726 1832 794
rect 420 480 1062 698
rect 1318 498 1832 726
rect 1320 482 1832 498
rect 420 420 926 480
rect 1484 452 1832 482
rect -1720 -366 -822 194
rect -1720 -582 -632 -366
rect -1720 -698 -768 -582
rect -1720 -2190 -1552 -698
rect -1274 -1402 -768 -698
rect -1720 -2358 -822 -2190
rect -1720 -2760 -1508 -2358
rect -990 -2760 -822 -2358
rect -1720 -2928 -822 -2760
<< pwell >>
rect -1508 3144 -990 3546
rect -1508 194 -990 596
rect -1508 -2760 -990 -2358
<< mvnmos >>
rect -1220 3850 -1120 4050
rect -932 3850 -832 3934
rect -1378 3262 -1278 3362
rect -1220 3262 -1120 3362
rect 1532 2016 1632 2216
rect 1690 2016 1790 2216
rect 2432 2016 2532 2216
rect 2590 2016 2690 2216
rect 3494 2006 3594 2206
rect 544 1500 644 1700
rect 702 1500 802 1700
rect 1532 1114 1632 1314
rect 1690 1114 1790 1314
rect -1220 900 -1120 1100
rect -932 900 -832 984
rect 2428 958 2528 1158
rect 2586 958 2686 1158
rect 3494 948 3594 1148
rect -1378 312 -1278 412
rect -1220 312 -1120 412
rect 544 152 644 352
rect 702 152 802 352
rect 1608 142 1708 342
rect -1220 -2054 -1120 -1854
rect -932 -2054 -832 -1970
rect -1378 -2642 -1278 -2542
rect -1220 -2642 -1120 -2542
<< mvpmos >>
rect -1596 5372 -1496 5472
rect -1438 5372 -1338 5472
rect -1150 4568 -1050 5468
rect -992 4568 -892 5468
rect -1596 2422 -1496 2522
rect -1438 2422 -1338 2522
rect -1150 1618 -1050 2518
rect -992 1618 -892 2518
rect 1532 2350 1632 2550
rect 1690 2350 1790 2550
rect 2432 2350 2532 2550
rect 2590 2350 2690 2550
rect 3494 2382 3594 2582
rect 544 1834 644 2034
rect 702 1834 802 2034
rect 1532 1448 1632 1648
rect 1690 1448 1790 1648
rect 2428 1292 2528 1492
rect 2586 1292 2686 1492
rect 3494 1324 3594 1524
rect 544 486 644 686
rect 702 486 802 686
rect 1608 518 1708 718
rect -1596 -532 -1496 -432
rect -1438 -532 -1338 -432
rect -1150 -1336 -1050 -436
rect -992 -1336 -892 -436
<< mvndiff >>
rect -1278 4038 -1220 4050
rect -1278 3862 -1266 4038
rect -1232 3862 -1220 4038
rect -1278 3850 -1220 3862
rect -1120 4038 -1062 4050
rect -1120 3862 -1108 4038
rect -1074 3862 -1062 4038
rect -1120 3850 -1062 3862
rect -990 3922 -932 3934
rect -990 3862 -978 3922
rect -944 3862 -932 3922
rect -990 3850 -932 3862
rect -832 3922 -774 3934
rect -832 3862 -820 3922
rect -786 3862 -774 3922
rect -832 3850 -774 3862
rect -1436 3350 -1378 3362
rect -1436 3274 -1424 3350
rect -1390 3274 -1378 3350
rect -1436 3262 -1378 3274
rect -1278 3350 -1220 3362
rect -1278 3274 -1266 3350
rect -1232 3274 -1220 3350
rect -1278 3262 -1220 3274
rect -1120 3350 -1062 3362
rect -1120 3274 -1108 3350
rect -1074 3274 -1062 3350
rect -1120 3262 -1062 3274
rect 1474 2204 1532 2216
rect 1474 2028 1486 2204
rect 1520 2028 1532 2204
rect 1474 2016 1532 2028
rect 1632 2204 1690 2216
rect 1632 2028 1644 2204
rect 1678 2028 1690 2204
rect 1632 2016 1690 2028
rect 1790 2204 1848 2216
rect 1790 2028 1802 2204
rect 1836 2028 1848 2204
rect 2374 2204 2432 2216
rect 1790 2016 1848 2028
rect 2374 2028 2386 2204
rect 2420 2028 2432 2204
rect 2374 2016 2432 2028
rect 2532 2204 2590 2216
rect 2532 2028 2544 2204
rect 2578 2028 2590 2204
rect 2532 2016 2590 2028
rect 2690 2204 2748 2216
rect 2690 2028 2702 2204
rect 2736 2028 2748 2204
rect 3436 2194 3494 2206
rect 2690 2016 2748 2028
rect 3436 2018 3448 2194
rect 3482 2018 3494 2194
rect 3436 2006 3494 2018
rect 3594 2194 3652 2206
rect 3594 2018 3606 2194
rect 3640 2018 3652 2194
rect 3594 2006 3652 2018
rect 486 1688 544 1700
rect 486 1512 498 1688
rect 532 1512 544 1688
rect 486 1500 544 1512
rect 644 1688 702 1700
rect 644 1512 656 1688
rect 690 1512 702 1688
rect 644 1500 702 1512
rect 802 1688 860 1700
rect 802 1512 814 1688
rect 848 1512 860 1688
rect 802 1500 860 1512
rect 1474 1302 1532 1314
rect 1474 1126 1486 1302
rect 1520 1126 1532 1302
rect 1474 1114 1532 1126
rect 1632 1302 1690 1314
rect 1632 1126 1644 1302
rect 1678 1126 1690 1302
rect 1632 1114 1690 1126
rect 1790 1302 1848 1314
rect 1790 1126 1802 1302
rect 1836 1126 1848 1302
rect 2370 1146 2428 1158
rect 1790 1114 1848 1126
rect -1278 1088 -1220 1100
rect -1278 912 -1266 1088
rect -1232 912 -1220 1088
rect -1278 900 -1220 912
rect -1120 1088 -1062 1100
rect -1120 912 -1108 1088
rect -1074 912 -1062 1088
rect -1120 900 -1062 912
rect -990 972 -932 984
rect -990 912 -978 972
rect -944 912 -932 972
rect -990 900 -932 912
rect -832 972 -774 984
rect -832 912 -820 972
rect -786 912 -774 972
rect 2370 970 2382 1146
rect 2416 970 2428 1146
rect 2370 958 2428 970
rect 2528 1146 2586 1158
rect 2528 970 2540 1146
rect 2574 970 2586 1146
rect 2528 958 2586 970
rect 2686 1146 2744 1158
rect 2686 970 2698 1146
rect 2732 970 2744 1146
rect 3436 1136 3494 1148
rect 2686 958 2744 970
rect 3436 960 3448 1136
rect 3482 960 3494 1136
rect -832 900 -774 912
rect 3436 948 3494 960
rect 3594 1136 3652 1148
rect 3594 960 3606 1136
rect 3640 960 3652 1136
rect 3594 948 3652 960
rect -1436 400 -1378 412
rect -1436 324 -1424 400
rect -1390 324 -1378 400
rect -1436 312 -1378 324
rect -1278 400 -1220 412
rect -1278 324 -1266 400
rect -1232 324 -1220 400
rect -1278 312 -1220 324
rect -1120 400 -1062 412
rect -1120 324 -1108 400
rect -1074 324 -1062 400
rect -1120 312 -1062 324
rect 486 340 544 352
rect 486 164 498 340
rect 532 164 544 340
rect 486 152 544 164
rect 644 340 702 352
rect 644 164 656 340
rect 690 164 702 340
rect 644 152 702 164
rect 802 340 860 352
rect 802 164 814 340
rect 848 164 860 340
rect 1550 330 1608 342
rect 802 152 860 164
rect 1550 154 1562 330
rect 1596 154 1608 330
rect 1550 142 1608 154
rect 1708 330 1766 342
rect 1708 154 1720 330
rect 1754 154 1766 330
rect 1708 142 1766 154
rect -1278 -1866 -1220 -1854
rect -1278 -2042 -1266 -1866
rect -1232 -2042 -1220 -1866
rect -1278 -2054 -1220 -2042
rect -1120 -1866 -1062 -1854
rect -1120 -2042 -1108 -1866
rect -1074 -2042 -1062 -1866
rect -1120 -2054 -1062 -2042
rect -990 -1982 -932 -1970
rect -990 -2042 -978 -1982
rect -944 -2042 -932 -1982
rect -990 -2054 -932 -2042
rect -832 -1982 -774 -1970
rect -832 -2042 -820 -1982
rect -786 -2042 -774 -1982
rect -832 -2054 -774 -2042
rect -1436 -2554 -1378 -2542
rect -1436 -2630 -1424 -2554
rect -1390 -2630 -1378 -2554
rect -1436 -2642 -1378 -2630
rect -1278 -2554 -1220 -2542
rect -1278 -2630 -1266 -2554
rect -1232 -2630 -1220 -2554
rect -1278 -2642 -1220 -2630
rect -1120 -2554 -1062 -2542
rect -1120 -2630 -1108 -2554
rect -1074 -2630 -1062 -2554
rect -1120 -2642 -1062 -2630
<< mvpdiff >>
rect -1654 5460 -1596 5472
rect -1654 5384 -1642 5460
rect -1608 5384 -1596 5460
rect -1654 5372 -1596 5384
rect -1496 5460 -1438 5472
rect -1496 5384 -1484 5460
rect -1450 5384 -1438 5460
rect -1496 5372 -1438 5384
rect -1338 5460 -1280 5472
rect -1338 5384 -1326 5460
rect -1292 5384 -1280 5460
rect -1338 5372 -1280 5384
rect -1208 5456 -1150 5468
rect -1208 4580 -1196 5456
rect -1162 4580 -1150 5456
rect -1208 4568 -1150 4580
rect -1050 5456 -992 5468
rect -1050 4580 -1038 5456
rect -1004 4580 -992 5456
rect -1050 4568 -992 4580
rect -892 5456 -834 5468
rect -892 4580 -880 5456
rect -846 4580 -834 5456
rect -892 4568 -834 4580
rect 3436 2570 3494 2582
rect -1654 2510 -1596 2522
rect -1654 2434 -1642 2510
rect -1608 2434 -1596 2510
rect -1654 2422 -1596 2434
rect -1496 2510 -1438 2522
rect -1496 2434 -1484 2510
rect -1450 2434 -1438 2510
rect -1496 2422 -1438 2434
rect -1338 2510 -1280 2522
rect 1474 2538 1532 2550
rect -1338 2434 -1326 2510
rect -1292 2434 -1280 2510
rect -1338 2422 -1280 2434
rect -1208 2506 -1150 2518
rect -1208 1630 -1196 2506
rect -1162 1630 -1150 2506
rect -1208 1618 -1150 1630
rect -1050 2506 -992 2518
rect -1050 1630 -1038 2506
rect -1004 1630 -992 2506
rect -1050 1618 -992 1630
rect -892 2506 -834 2518
rect -892 1630 -880 2506
rect -846 1630 -834 2506
rect 1474 2362 1486 2538
rect 1520 2362 1532 2538
rect 1474 2350 1532 2362
rect 1632 2538 1690 2550
rect 1632 2362 1644 2538
rect 1678 2362 1690 2538
rect 1632 2350 1690 2362
rect 1790 2538 1848 2550
rect 1790 2362 1802 2538
rect 1836 2362 1848 2538
rect 2374 2538 2432 2550
rect 1790 2350 1848 2362
rect 2374 2362 2386 2538
rect 2420 2362 2432 2538
rect 2374 2350 2432 2362
rect 2532 2538 2590 2550
rect 2532 2362 2544 2538
rect 2578 2362 2590 2538
rect 2532 2350 2590 2362
rect 2690 2538 2748 2550
rect 2690 2362 2702 2538
rect 2736 2362 2748 2538
rect 3436 2394 3448 2570
rect 3482 2394 3494 2570
rect 3436 2382 3494 2394
rect 3594 2570 3652 2582
rect 3594 2394 3606 2570
rect 3640 2394 3652 2570
rect 3594 2382 3652 2394
rect 2690 2350 2748 2362
rect 486 2022 544 2034
rect 486 1846 498 2022
rect 532 1846 544 2022
rect 486 1834 544 1846
rect 644 2022 702 2034
rect 644 1846 656 2022
rect 690 1846 702 2022
rect 644 1834 702 1846
rect 802 2022 860 2034
rect 802 1846 814 2022
rect 848 1846 860 2022
rect 802 1834 860 1846
rect -892 1618 -834 1630
rect 1474 1636 1532 1648
rect 1474 1460 1486 1636
rect 1520 1460 1532 1636
rect 1474 1448 1532 1460
rect 1632 1636 1690 1648
rect 1632 1460 1644 1636
rect 1678 1460 1690 1636
rect 1632 1448 1690 1460
rect 1790 1636 1848 1648
rect 1790 1460 1802 1636
rect 1836 1460 1848 1636
rect 3436 1512 3494 1524
rect 1790 1448 1848 1460
rect 2370 1480 2428 1492
rect 2370 1304 2382 1480
rect 2416 1304 2428 1480
rect 2370 1292 2428 1304
rect 2528 1480 2586 1492
rect 2528 1304 2540 1480
rect 2574 1304 2586 1480
rect 2528 1292 2586 1304
rect 2686 1480 2744 1492
rect 2686 1304 2698 1480
rect 2732 1304 2744 1480
rect 3436 1336 3448 1512
rect 3482 1336 3494 1512
rect 3436 1324 3494 1336
rect 3594 1512 3652 1524
rect 3594 1336 3606 1512
rect 3640 1336 3652 1512
rect 3594 1324 3652 1336
rect 2686 1292 2744 1304
rect 1550 706 1608 718
rect 486 674 544 686
rect 486 498 498 674
rect 532 498 544 674
rect 486 486 544 498
rect 644 674 702 686
rect 644 498 656 674
rect 690 498 702 674
rect 644 486 702 498
rect 802 674 860 686
rect 802 498 814 674
rect 848 498 860 674
rect 1550 530 1562 706
rect 1596 530 1608 706
rect 1550 518 1608 530
rect 1708 706 1766 718
rect 1708 530 1720 706
rect 1754 530 1766 706
rect 1708 518 1766 530
rect 802 486 860 498
rect -1654 -444 -1596 -432
rect -1654 -520 -1642 -444
rect -1608 -520 -1596 -444
rect -1654 -532 -1596 -520
rect -1496 -444 -1438 -432
rect -1496 -520 -1484 -444
rect -1450 -520 -1438 -444
rect -1496 -532 -1438 -520
rect -1338 -444 -1280 -432
rect -1338 -520 -1326 -444
rect -1292 -520 -1280 -444
rect -1338 -532 -1280 -520
rect -1208 -448 -1150 -436
rect -1208 -1324 -1196 -448
rect -1162 -1324 -1150 -448
rect -1208 -1336 -1150 -1324
rect -1050 -448 -992 -436
rect -1050 -1324 -1038 -448
rect -1004 -1324 -992 -448
rect -1050 -1336 -992 -1324
rect -892 -448 -834 -436
rect -892 -1324 -880 -448
rect -846 -1324 -834 -448
rect -892 -1336 -834 -1324
<< mvndiffc >>
rect -1266 3862 -1232 4038
rect -1108 3862 -1074 4038
rect -978 3862 -944 3922
rect -820 3862 -786 3922
rect -1424 3274 -1390 3350
rect -1266 3274 -1232 3350
rect -1108 3274 -1074 3350
rect 1486 2028 1520 2204
rect 1644 2028 1678 2204
rect 1802 2028 1836 2204
rect 2386 2028 2420 2204
rect 2544 2028 2578 2204
rect 2702 2028 2736 2204
rect 3448 2018 3482 2194
rect 3606 2018 3640 2194
rect 498 1512 532 1688
rect 656 1512 690 1688
rect 814 1512 848 1688
rect 1486 1126 1520 1302
rect 1644 1126 1678 1302
rect 1802 1126 1836 1302
rect -1266 912 -1232 1088
rect -1108 912 -1074 1088
rect -978 912 -944 972
rect -820 912 -786 972
rect 2382 970 2416 1146
rect 2540 970 2574 1146
rect 2698 970 2732 1146
rect 3448 960 3482 1136
rect 3606 960 3640 1136
rect -1424 324 -1390 400
rect -1266 324 -1232 400
rect -1108 324 -1074 400
rect 498 164 532 340
rect 656 164 690 340
rect 814 164 848 340
rect 1562 154 1596 330
rect 1720 154 1754 330
rect -1266 -2042 -1232 -1866
rect -1108 -2042 -1074 -1866
rect -978 -2042 -944 -1982
rect -820 -2042 -786 -1982
rect -1424 -2630 -1390 -2554
rect -1266 -2630 -1232 -2554
rect -1108 -2630 -1074 -2554
<< mvpdiffc >>
rect -1642 5384 -1608 5460
rect -1484 5384 -1450 5460
rect -1326 5384 -1292 5460
rect -1196 4580 -1162 5456
rect -1038 4580 -1004 5456
rect -880 4580 -846 5456
rect -1642 2434 -1608 2510
rect -1484 2434 -1450 2510
rect -1326 2434 -1292 2510
rect -1196 1630 -1162 2506
rect -1038 1630 -1004 2506
rect -880 1630 -846 2506
rect 1486 2362 1520 2538
rect 1644 2362 1678 2538
rect 1802 2362 1836 2538
rect 2386 2362 2420 2538
rect 2544 2362 2578 2538
rect 2702 2362 2736 2538
rect 3448 2394 3482 2570
rect 3606 2394 3640 2570
rect 498 1846 532 2022
rect 656 1846 690 2022
rect 814 1846 848 2022
rect 1486 1460 1520 1636
rect 1644 1460 1678 1636
rect 1802 1460 1836 1636
rect 2382 1304 2416 1480
rect 2540 1304 2574 1480
rect 2698 1304 2732 1480
rect 3448 1336 3482 1512
rect 3606 1336 3640 1512
rect 498 498 532 674
rect 656 498 690 674
rect 814 498 848 674
rect 1562 530 1596 706
rect 1720 530 1754 706
rect -1642 -520 -1608 -444
rect -1484 -520 -1450 -444
rect -1326 -520 -1292 -444
rect -1196 -1324 -1162 -448
rect -1038 -1324 -1004 -448
rect -880 -1324 -846 -448
<< mvpsubdiff >>
rect -1132 4172 -1050 4182
rect -1132 4134 -1108 4172
rect -1074 4134 -1050 4172
rect -1132 4124 -1050 4134
rect -1290 3512 -1208 3520
rect -1290 3442 -1266 3512
rect -1232 3442 -1208 3512
rect -1290 3436 -1208 3442
rect -2626 2160 -2534 2180
rect -2626 2076 -2602 2160
rect -2558 2076 -2534 2160
rect -2626 2056 -2534 2076
rect 1922 2112 2004 2126
rect 1922 2054 1946 2112
rect 1980 2054 2004 2112
rect 1922 2040 2004 2054
rect 3198 2152 3338 2192
rect 2822 2112 2904 2126
rect 2822 2054 2846 2112
rect 2880 2054 2904 2112
rect 2822 2040 2904 2054
rect 3198 2072 3238 2152
rect 3298 2072 3338 2152
rect 3198 2032 3338 2072
rect 934 1596 1016 1610
rect 934 1538 958 1596
rect 992 1538 1016 1596
rect 934 1524 1016 1538
rect -1132 1222 -1050 1232
rect -1132 1184 -1108 1222
rect -1074 1184 -1050 1222
rect -1132 1174 -1050 1184
rect 1922 1210 2004 1224
rect 1922 1152 1946 1210
rect 1980 1152 2004 1210
rect 1922 1138 2004 1152
rect 3198 1094 3338 1134
rect 2818 1054 2900 1068
rect 2818 996 2842 1054
rect 2876 996 2900 1054
rect 2818 982 2900 996
rect 3198 1014 3238 1094
rect 3298 1014 3338 1094
rect 3198 974 3338 1014
rect -2626 694 -2534 718
rect -2626 610 -2602 694
rect -2558 610 -2534 694
rect -2626 586 -2534 610
rect -1290 562 -1208 570
rect -1290 492 -1266 562
rect -1232 492 -1208 562
rect -1290 486 -1208 492
rect 1312 288 1452 328
rect 934 248 1016 262
rect 934 190 958 248
rect 992 190 1016 248
rect 934 176 1016 190
rect 1312 208 1352 288
rect 1412 208 1452 288
rect 1312 168 1452 208
rect -2626 -774 -2534 -750
rect -2626 -858 -2602 -774
rect -2558 -858 -2534 -774
rect -2626 -882 -2534 -858
rect -1132 -1732 -1050 -1722
rect -1132 -1770 -1108 -1732
rect -1074 -1770 -1050 -1732
rect -1132 -1780 -1050 -1770
rect -2412 -2120 -2320 -2096
rect -2412 -2204 -2388 -2120
rect -2344 -2204 -2320 -2120
rect -2412 -2228 -2320 -2204
rect -1290 -2392 -1208 -2384
rect -1290 -2462 -1266 -2392
rect -1232 -2462 -1208 -2392
rect -1290 -2468 -1208 -2462
<< mvnsubdiff >>
rect -780 5448 -698 5472
rect -780 5412 -756 5448
rect -722 5412 -698 5448
rect -780 5388 -698 5412
rect -780 2498 -698 2522
rect -780 2462 -756 2498
rect -722 2462 -698 2498
rect -780 2438 -698 2462
rect 1902 2482 1984 2496
rect 1902 2424 1926 2482
rect 1960 2424 1984 2482
rect 1902 2410 1984 2424
rect 3272 2508 3354 2522
rect 2802 2482 2884 2496
rect 2802 2424 2826 2482
rect 2860 2424 2884 2482
rect 2802 2410 2884 2424
rect 3272 2436 3296 2508
rect 3330 2436 3354 2508
rect 3272 2412 3354 2436
rect 914 1966 996 1980
rect 914 1908 938 1966
rect 972 1908 996 1966
rect 914 1894 996 1908
rect 1902 1580 1984 1594
rect 1902 1522 1926 1580
rect 1960 1522 1984 1580
rect 1902 1508 1984 1522
rect 3272 1450 3354 1464
rect 2798 1424 2880 1438
rect 2798 1366 2822 1424
rect 2856 1366 2880 1424
rect 2798 1352 2880 1366
rect 3272 1378 3296 1450
rect 3330 1378 3354 1450
rect 3272 1354 3354 1378
rect 1386 644 1468 658
rect 914 618 996 632
rect 914 560 938 618
rect 972 560 996 618
rect 914 546 996 560
rect 1386 572 1410 644
rect 1444 572 1468 644
rect 1386 548 1468 572
rect -780 -456 -698 -432
rect -780 -492 -756 -456
rect -722 -492 -698 -456
rect -780 -516 -698 -492
<< mvpsubdiffcont >>
rect -1108 4134 -1074 4172
rect -1266 3442 -1232 3512
rect -2602 2076 -2558 2160
rect 1946 2054 1980 2112
rect 2846 2054 2880 2112
rect 3238 2072 3298 2152
rect 958 1538 992 1596
rect -1108 1184 -1074 1222
rect 1946 1152 1980 1210
rect 2842 996 2876 1054
rect 3238 1014 3298 1094
rect -2602 610 -2558 694
rect -1266 492 -1232 562
rect 958 190 992 248
rect 1352 208 1412 288
rect -2602 -858 -2558 -774
rect -1108 -1770 -1074 -1732
rect -2388 -2204 -2344 -2120
rect -1266 -2462 -1232 -2392
<< mvnsubdiffcont >>
rect -756 5412 -722 5448
rect -756 2462 -722 2498
rect 1926 2424 1960 2482
rect 2826 2424 2860 2482
rect 3296 2436 3330 2508
rect 938 1908 972 1966
rect 1926 1522 1960 1580
rect 2822 1366 2856 1424
rect 3296 1378 3330 1450
rect 938 560 972 618
rect 1410 572 1444 644
rect -756 -492 -722 -456
<< poly >>
rect -1596 5472 -1496 5498
rect -1438 5472 -1338 5498
rect -1150 5468 -1050 5494
rect -992 5468 -892 5494
rect -1596 5346 -1496 5372
rect -1438 5346 -1338 5372
rect -1654 5322 -1338 5346
rect -1654 5284 -1642 5322
rect -1608 5284 -1428 5322
rect -1654 5282 -1428 5284
rect -1388 5282 -1338 5322
rect -1654 5258 -1338 5282
rect -1150 4546 -1050 4568
rect -992 4546 -892 4568
rect -1208 4518 -892 4546
rect -1208 4484 -1174 4518
rect -1128 4484 -892 4518
rect -1208 4458 -892 4484
rect -1220 4050 -1120 4076
rect -932 3934 -832 3960
rect -1220 3824 -1120 3850
rect -932 3824 -832 3850
rect -1220 3802 -832 3824
rect -1220 3766 -882 3802
rect -844 3766 -832 3802
rect -1220 3742 -832 3766
rect -1080 3692 -980 3742
rect -1378 3362 -1278 3388
rect -1220 3362 -1120 3388
rect -1378 3160 -1278 3262
rect -1378 3124 -1346 3160
rect -1308 3124 -1278 3160
rect -1378 3102 -1278 3124
rect -1220 3156 -1120 3262
rect -1220 3120 -1190 3156
rect -1152 3120 -1120 3156
rect -1220 3102 -1120 3120
rect 3494 2582 3594 2608
rect 1532 2550 1632 2576
rect 1690 2550 1790 2576
rect 2432 2550 2532 2576
rect 2590 2550 2690 2576
rect -1596 2522 -1496 2548
rect -1438 2522 -1338 2548
rect -1150 2518 -1050 2544
rect -992 2518 -892 2544
rect -1596 2396 -1496 2422
rect -1438 2396 -1338 2422
rect -1654 2372 -1338 2396
rect -1654 2334 -1642 2372
rect -1608 2334 -1428 2372
rect -1654 2332 -1428 2334
rect -1388 2332 -1338 2372
rect -1654 2308 -1338 2332
rect 1532 2216 1632 2350
rect 1690 2216 1790 2350
rect 2432 2216 2532 2350
rect 2590 2216 2690 2350
rect 3494 2304 3594 2382
rect 3494 2270 3522 2304
rect 3558 2270 3594 2304
rect 544 2034 644 2060
rect 702 2034 802 2060
rect 3494 2206 3594 2270
rect 1532 1978 1632 2016
rect 1532 1944 1562 1978
rect 1598 1944 1632 1978
rect 1532 1934 1632 1944
rect 1690 1978 1790 2016
rect 1690 1944 1718 1978
rect 1754 1944 1790 1978
rect 1690 1934 1790 1944
rect 2432 1978 2532 2016
rect 2432 1944 2462 1978
rect 2498 1944 2532 1978
rect 2432 1934 2532 1944
rect 2590 1978 2690 2016
rect 3494 1980 3594 2006
rect 2590 1944 2618 1978
rect 2654 1944 2690 1978
rect 2590 1934 2690 1944
rect 544 1700 644 1834
rect 702 1700 802 1834
rect -1150 1596 -1050 1618
rect -992 1596 -892 1618
rect -1208 1568 -892 1596
rect -1208 1534 -1174 1568
rect -1128 1534 -892 1568
rect -1208 1508 -892 1534
rect 1532 1648 1632 1674
rect 1690 1648 1790 1674
rect 544 1462 644 1500
rect 544 1428 576 1462
rect 612 1428 644 1462
rect 544 1418 644 1428
rect 702 1462 802 1500
rect 702 1428 730 1462
rect 766 1428 802 1462
rect 3494 1524 3594 1550
rect 2428 1492 2528 1518
rect 2586 1492 2686 1518
rect 702 1418 802 1428
rect 1532 1314 1632 1448
rect 1690 1314 1790 1448
rect -1220 1100 -1120 1126
rect 2428 1158 2528 1292
rect 2586 1158 2686 1292
rect 3494 1246 3594 1324
rect 3494 1212 3522 1246
rect 3558 1212 3594 1246
rect 1532 1076 1632 1114
rect 1532 1042 1562 1076
rect 1598 1042 1632 1076
rect 1532 1032 1632 1042
rect 1690 1076 1790 1114
rect 1690 1042 1718 1076
rect 1754 1042 1790 1076
rect 1690 1032 1790 1042
rect -932 984 -832 1010
rect 3494 1148 3594 1212
rect 2428 920 2528 958
rect -1220 874 -1120 900
rect -932 874 -832 900
rect 2428 886 2458 920
rect 2494 886 2528 920
rect 2428 876 2528 886
rect 2586 920 2686 958
rect 3494 922 3594 948
rect 2586 886 2614 920
rect 2650 886 2686 920
rect 2586 876 2686 886
rect -1220 854 -832 874
rect -1220 818 -900 854
rect -862 818 -832 854
rect -1220 792 -832 818
rect -1080 742 -980 792
rect 1608 718 1708 744
rect 544 686 644 712
rect 702 686 802 712
rect -1378 412 -1278 438
rect -1220 412 -1120 438
rect 544 352 644 486
rect 702 352 802 486
rect 1608 440 1708 518
rect 1608 406 1636 440
rect 1672 406 1708 440
rect -1378 210 -1278 312
rect -1378 174 -1346 210
rect -1308 174 -1278 210
rect -1378 152 -1278 174
rect -1220 206 -1120 312
rect -1220 172 -1188 206
rect -1150 172 -1120 206
rect -1220 152 -1120 172
rect 1608 342 1708 406
rect 544 114 644 152
rect 544 80 574 114
rect 610 80 644 114
rect 544 70 644 80
rect 702 114 802 152
rect 1608 116 1708 142
rect 702 80 730 114
rect 766 80 802 114
rect 702 70 802 80
rect -1596 -432 -1496 -406
rect -1438 -432 -1338 -406
rect -1150 -436 -1050 -410
rect -992 -436 -892 -410
rect -1596 -558 -1496 -532
rect -1438 -558 -1338 -532
rect -1654 -582 -1338 -558
rect -1654 -620 -1642 -582
rect -1608 -620 -1428 -582
rect -1654 -622 -1428 -620
rect -1388 -622 -1338 -582
rect -1654 -646 -1338 -622
rect -1150 -1358 -1050 -1336
rect -992 -1358 -892 -1336
rect -1208 -1386 -892 -1358
rect -1208 -1420 -1174 -1386
rect -1128 -1420 -892 -1386
rect -1208 -1446 -892 -1420
rect -1220 -1854 -1120 -1828
rect -932 -1970 -832 -1944
rect -1220 -2080 -1120 -2054
rect -932 -2080 -832 -2054
rect -1220 -2124 -832 -2080
rect -1220 -2160 -1048 -2124
rect -1010 -2160 -832 -2124
rect -1220 -2162 -832 -2160
rect -1080 -2212 -980 -2162
rect -1378 -2542 -1278 -2516
rect -1220 -2542 -1120 -2516
rect -1378 -2746 -1278 -2642
rect -1378 -2782 -1348 -2746
rect -1310 -2782 -1278 -2746
rect -1378 -2802 -1278 -2782
rect -1220 -2748 -1120 -2642
rect -1220 -2784 -1190 -2748
rect -1152 -2784 -1120 -2748
rect -1220 -2802 -1120 -2784
<< polycont >>
rect -1642 5284 -1608 5322
rect -1428 5282 -1388 5322
rect -1174 4484 -1128 4518
rect -882 3766 -844 3802
rect -1346 3124 -1308 3160
rect -1190 3120 -1152 3156
rect -1642 2334 -1608 2372
rect -1428 2332 -1388 2372
rect 3522 2270 3558 2304
rect 1562 1944 1598 1978
rect 1718 1944 1754 1978
rect 2462 1944 2498 1978
rect 2618 1944 2654 1978
rect -1174 1534 -1128 1568
rect 576 1428 612 1462
rect 730 1428 766 1462
rect 3522 1212 3558 1246
rect 1562 1042 1598 1076
rect 1718 1042 1754 1076
rect 2458 886 2494 920
rect 2614 886 2650 920
rect -900 818 -862 854
rect 1636 406 1672 440
rect -1346 174 -1308 210
rect -1188 172 -1150 206
rect 574 80 610 114
rect 730 80 766 114
rect -1642 -620 -1608 -582
rect -1428 -622 -1388 -582
rect -1174 -1420 -1128 -1386
rect -1048 -2160 -1010 -2124
rect -1348 -2782 -1310 -2746
rect -1190 -2784 -1152 -2748
<< xpolycontact >>
rect -2474 2818 -1904 3250
rect -2474 2282 -1904 2714
rect -2474 1530 -1904 1962
rect -2474 850 -1904 1282
rect -2476 34 -1906 466
rect -2476 -646 -1906 -214
rect -2476 -1406 -1906 -974
rect -2476 -1942 -1906 -1510
<< xpolyres >>
rect -2474 2714 -1904 2818
rect -2474 1282 -1904 1530
rect -2476 -214 -1906 34
rect -2476 -1510 -1906 -1406
<< locali >>
rect -1642 5460 -1608 5476
rect -1642 5322 -1608 5384
rect -1484 5460 -1450 5476
rect -1484 5368 -1450 5384
rect -1326 5460 -1292 5476
rect -1326 5368 -1292 5384
rect -1196 5456 -1162 5472
rect -1642 5268 -1608 5284
rect -1428 5322 -1388 5338
rect -1428 5266 -1388 5282
rect -1196 4564 -1162 4580
rect -1038 5456 -1004 5472
rect -1038 4564 -1004 4580
rect -880 5456 -846 5472
rect -756 5448 -722 5468
rect -846 5412 -756 5448
rect -756 5392 -722 5412
rect -880 4564 -846 4580
rect -1328 4530 -1288 4542
rect -1328 4478 -1288 4490
rect -1190 4484 -1174 4518
rect -1128 4484 -1112 4518
rect -1108 4172 -1074 4196
rect -1266 4038 -1232 4054
rect -1266 3846 -1232 3862
rect -1108 4038 -1074 4134
rect -1108 3846 -1074 3862
rect -978 3922 -944 3938
rect -978 3846 -944 3862
rect -820 3922 -786 3938
rect -820 3846 -786 3862
rect -882 3802 -844 3818
rect -882 3750 -844 3766
rect -1266 3512 -1232 3528
rect -1424 3350 -1390 3366
rect -1424 3258 -1390 3274
rect -1266 3350 -1232 3442
rect -1266 3258 -1232 3274
rect -1108 3350 -1074 3366
rect -1108 3258 -1074 3274
rect -1346 3160 -1308 3176
rect -1346 3104 -1308 3124
rect -1190 3156 -1152 3172
rect -1190 3104 -1152 3120
rect 3448 2570 3482 2586
rect 1486 2538 1520 2554
rect -1642 2510 -1608 2526
rect -1642 2372 -1608 2434
rect -1484 2510 -1450 2526
rect -1484 2418 -1450 2434
rect -1326 2510 -1292 2526
rect -1326 2418 -1292 2434
rect -1196 2506 -1162 2522
rect -1642 2318 -1608 2334
rect -1428 2372 -1388 2388
rect -1428 2316 -1388 2332
rect -2602 2160 -2558 2180
rect -2602 2056 -2558 2076
rect -1196 1614 -1162 1630
rect -1038 2506 -1004 2522
rect -1038 1614 -1004 1630
rect -880 2506 -846 2522
rect -756 2498 -722 2518
rect -846 2462 -756 2498
rect -756 2442 -722 2462
rect 1486 2346 1520 2362
rect 1644 2538 1678 2554
rect 1644 2346 1678 2362
rect 1802 2538 1836 2554
rect 2386 2538 2420 2554
rect 1926 2482 1960 2500
rect 1836 2432 1926 2470
rect 1926 2406 1960 2424
rect 1802 2346 1836 2362
rect 2386 2346 2420 2362
rect 2544 2538 2578 2554
rect 2544 2346 2578 2362
rect 2702 2538 2736 2554
rect 3296 2508 3330 2536
rect 2826 2482 2860 2500
rect 2736 2432 2826 2470
rect 2826 2406 2860 2424
rect 3330 2452 3448 2498
rect 3296 2410 3330 2436
rect 3448 2378 3482 2394
rect 3606 2570 3640 2586
rect 3606 2378 3640 2394
rect 2702 2346 2736 2362
rect 3522 2304 3558 2320
rect 3522 2252 3558 2270
rect 1486 2204 1520 2220
rect 498 2022 532 2038
rect 498 1830 532 1846
rect 656 2022 690 2038
rect 656 1830 690 1846
rect 814 2022 848 2038
rect 1486 2012 1520 2028
rect 1644 2204 1678 2220
rect 1644 2012 1678 2028
rect 1802 2204 1836 2220
rect 2386 2204 2420 2220
rect 1946 2112 1980 2136
rect 1836 2062 1946 2100
rect 1946 2030 1980 2054
rect 1802 2012 1836 2028
rect 2386 2012 2420 2028
rect 2544 2204 2578 2220
rect 2544 2012 2578 2028
rect 2702 2204 2736 2220
rect 3448 2194 3482 2210
rect 3218 2152 3318 2172
rect 2846 2112 2880 2136
rect 2736 2062 2846 2100
rect 2846 2030 2880 2054
rect 3218 2072 3238 2152
rect 3298 2072 3448 2152
rect 3218 2052 3318 2072
rect 2702 2012 2736 2028
rect 3448 2002 3482 2018
rect 3606 2194 3640 2210
rect 3606 2002 3640 2018
rect 938 1966 972 1984
rect 848 1916 938 1954
rect 1562 1978 1598 1994
rect 1562 1926 1598 1944
rect 1718 1978 1754 1994
rect 1718 1926 1754 1944
rect 2462 1978 2498 1994
rect 2462 1926 2498 1944
rect 2618 1978 2654 1994
rect 2618 1926 2654 1944
rect 938 1890 972 1908
rect 814 1830 848 1846
rect -880 1614 -846 1630
rect 498 1688 532 1704
rect -1328 1580 -1288 1592
rect -1328 1528 -1288 1540
rect -1190 1534 -1174 1568
rect -1128 1534 -1112 1568
rect 498 1496 532 1512
rect 656 1688 690 1704
rect 656 1496 690 1512
rect 814 1688 848 1704
rect 1486 1636 1520 1652
rect 958 1596 992 1620
rect 848 1546 958 1584
rect 958 1514 992 1538
rect 814 1496 848 1512
rect 576 1462 612 1478
rect 576 1410 612 1428
rect 730 1462 766 1478
rect 1486 1444 1520 1460
rect 1644 1636 1678 1652
rect 1644 1444 1678 1460
rect 1802 1636 1836 1652
rect 1926 1580 1960 1598
rect 1836 1530 1926 1568
rect 1926 1504 1960 1522
rect 3448 1512 3482 1528
rect 1802 1444 1836 1460
rect 2382 1480 2416 1496
rect 730 1410 766 1428
rect 1486 1302 1520 1318
rect -1108 1222 -1074 1246
rect -1266 1088 -1232 1104
rect -1266 896 -1232 912
rect -1108 1088 -1074 1184
rect 1486 1110 1520 1126
rect 1644 1302 1678 1318
rect 1644 1110 1678 1126
rect 1802 1302 1836 1318
rect 2382 1288 2416 1304
rect 2540 1480 2574 1496
rect 2540 1288 2574 1304
rect 2698 1480 2732 1496
rect 3296 1450 3330 1478
rect 2822 1424 2856 1442
rect 2732 1374 2822 1412
rect 2822 1348 2856 1366
rect 3330 1394 3448 1440
rect 3296 1352 3330 1378
rect 3448 1320 3482 1336
rect 3606 1512 3640 1528
rect 3606 1320 3640 1336
rect 2698 1288 2732 1304
rect 3522 1246 3558 1262
rect 1946 1210 1980 1234
rect 1836 1160 1946 1198
rect 3522 1194 3558 1212
rect 1946 1128 1980 1152
rect 2382 1146 2416 1162
rect 1802 1110 1836 1126
rect 1562 1076 1598 1092
rect 1562 1024 1598 1042
rect 1718 1076 1754 1092
rect 1718 1024 1754 1042
rect -1108 896 -1074 912
rect -978 972 -944 988
rect -978 896 -944 912
rect -820 972 -786 988
rect 2382 954 2416 970
rect 2540 1146 2574 1162
rect 2540 954 2574 970
rect 2698 1146 2732 1162
rect 3448 1136 3482 1152
rect 3218 1094 3318 1114
rect 2842 1054 2876 1078
rect 2732 1004 2842 1042
rect 2842 972 2876 996
rect 3218 1014 3238 1094
rect 3298 1014 3448 1094
rect 3218 994 3318 1014
rect 2698 954 2732 970
rect 3448 944 3482 960
rect 3606 1136 3640 1152
rect 3606 944 3640 960
rect -820 896 -786 912
rect 2458 920 2494 936
rect -900 854 -862 870
rect 2458 868 2494 886
rect 2614 920 2650 936
rect 2614 868 2650 886
rect -900 802 -862 818
rect -2602 694 -2558 718
rect 1562 706 1596 722
rect -2602 586 -2558 610
rect 498 674 532 690
rect -1266 562 -1232 578
rect -1424 400 -1390 416
rect -1424 308 -1390 324
rect -1266 400 -1232 492
rect 498 482 532 498
rect 656 674 690 690
rect 656 482 690 498
rect 814 674 848 690
rect 1410 644 1444 672
rect 938 618 972 636
rect 848 568 938 606
rect 938 542 972 560
rect 1444 588 1562 634
rect 1410 546 1444 572
rect 1562 514 1596 530
rect 1720 706 1754 722
rect 1720 514 1754 530
rect 814 482 848 498
rect 1636 440 1672 456
rect -1266 308 -1232 324
rect -1108 400 -1074 416
rect 1636 388 1672 406
rect -1108 308 -1074 324
rect 498 340 532 356
rect -1346 210 -1308 226
rect -1346 154 -1308 174
rect -1188 206 -1150 224
rect -1188 152 -1150 172
rect 498 148 532 164
rect 656 340 690 356
rect 656 148 690 164
rect 814 340 848 356
rect 1562 330 1596 346
rect 1332 288 1432 308
rect 958 248 992 272
rect 848 198 958 236
rect 958 166 992 190
rect 1332 208 1352 288
rect 1412 208 1562 288
rect 1332 188 1432 208
rect 814 148 848 164
rect 1562 138 1596 154
rect 1720 330 1754 346
rect 1720 138 1754 154
rect 574 114 610 130
rect 574 62 610 80
rect 730 114 766 130
rect 730 62 766 80
rect -1642 -444 -1608 -428
rect -1642 -582 -1608 -520
rect -1484 -444 -1450 -428
rect -1484 -536 -1450 -520
rect -1326 -444 -1292 -428
rect -1326 -536 -1292 -520
rect -1196 -448 -1162 -432
rect -1642 -636 -1608 -620
rect -1428 -582 -1388 -566
rect -1428 -638 -1388 -622
rect -2602 -774 -2558 -750
rect -2602 -882 -2558 -858
rect -1196 -1340 -1162 -1324
rect -1038 -448 -1004 -432
rect -1038 -1340 -1004 -1324
rect -880 -448 -846 -432
rect -756 -456 -722 -436
rect -846 -492 -756 -456
rect -756 -512 -722 -492
rect -880 -1340 -846 -1324
rect -1328 -1374 -1288 -1362
rect -1328 -1426 -1288 -1414
rect -1190 -1420 -1174 -1386
rect -1128 -1420 -1112 -1386
rect -1108 -1732 -1074 -1708
rect -1266 -1866 -1232 -1850
rect -1266 -2058 -1232 -2042
rect -1108 -1866 -1074 -1770
rect -1108 -2058 -1074 -2042
rect -978 -1982 -944 -1966
rect -978 -2058 -944 -2042
rect -820 -1982 -786 -1966
rect -820 -2058 -786 -2042
rect -2388 -2120 -2344 -2096
rect -1048 -2124 -1010 -2108
rect -1048 -2176 -1010 -2160
rect -2388 -2228 -2344 -2204
rect -1266 -2392 -1232 -2376
rect -1424 -2554 -1390 -2538
rect -1424 -2646 -1390 -2630
rect -1266 -2554 -1232 -2462
rect -1266 -2646 -1232 -2630
rect -1108 -2554 -1074 -2538
rect -1108 -2646 -1074 -2630
rect -1348 -2746 -1310 -2730
rect -1348 -2798 -1310 -2782
rect -1190 -2748 -1152 -2732
rect -1190 -2800 -1152 -2784
<< viali >>
rect -1642 5384 -1608 5460
rect -1484 5384 -1450 5460
rect -1326 5384 -1292 5460
rect -1428 5282 -1388 5322
rect -1196 4580 -1162 5456
rect -1038 4580 -1004 5456
rect -880 4580 -846 5456
rect -1328 4490 -1288 4530
rect -1174 4484 -1128 4518
rect -1266 3862 -1232 4038
rect -1108 3862 -1074 4038
rect -978 3862 -944 3922
rect -820 3862 -786 3922
rect -882 3766 -844 3802
rect -1424 3274 -1390 3350
rect -1266 3274 -1232 3350
rect -1108 3274 -1074 3350
rect -2458 2835 -1920 3232
rect -1346 3124 -1308 3160
rect -1190 3120 -1152 3156
rect -2458 2300 -1920 2697
rect -1642 2434 -1608 2510
rect -1484 2434 -1450 2510
rect -1326 2434 -1292 2510
rect -1428 2332 -1388 2372
rect -2602 2076 -2558 2160
rect -2458 1547 -1920 1944
rect -1196 1630 -1162 2506
rect -1038 1630 -1004 2506
rect -880 1630 -846 2506
rect 1486 2362 1520 2538
rect 1644 2362 1678 2538
rect 1802 2362 1836 2538
rect 2386 2362 2420 2538
rect 2544 2362 2578 2538
rect 2702 2362 2736 2538
rect 3448 2394 3482 2570
rect 3606 2394 3640 2570
rect 3522 2270 3558 2304
rect 498 1846 532 2022
rect 656 1846 690 2022
rect 814 1846 848 2022
rect 1486 2028 1520 2204
rect 1644 2028 1678 2204
rect 1802 2028 1836 2204
rect 2386 2028 2420 2204
rect 2544 2028 2578 2204
rect 2702 2028 2736 2204
rect 3448 2018 3482 2194
rect 3606 2018 3640 2194
rect 1562 1944 1598 1978
rect 1718 1944 1754 1978
rect 2462 1944 2498 1978
rect 2618 1944 2654 1978
rect -1328 1540 -1288 1580
rect -1174 1534 -1128 1568
rect 498 1512 532 1688
rect 656 1512 690 1688
rect 814 1512 848 1688
rect 576 1428 612 1462
rect 730 1428 766 1462
rect 1486 1460 1520 1636
rect 1644 1460 1678 1636
rect 1802 1460 1836 1636
rect -2458 868 -1920 1265
rect -1266 912 -1232 1088
rect 1486 1126 1520 1302
rect 1644 1126 1678 1302
rect 1802 1126 1836 1302
rect 2382 1304 2416 1480
rect 2540 1304 2574 1480
rect 2698 1304 2732 1480
rect 3448 1336 3482 1512
rect 3606 1336 3640 1512
rect 3522 1212 3558 1246
rect -1108 912 -1074 1088
rect 1562 1042 1598 1076
rect 1718 1042 1754 1076
rect -978 912 -944 972
rect -820 912 -786 972
rect 2382 970 2416 1146
rect 2540 970 2574 1146
rect 2698 970 2732 1146
rect 3448 960 3482 1136
rect 3606 960 3640 1136
rect 2458 886 2494 920
rect 2614 886 2650 920
rect -900 818 -862 854
rect -2602 610 -2558 694
rect -2460 51 -1922 448
rect -1424 324 -1390 400
rect 498 498 532 674
rect 656 498 690 674
rect 814 498 848 674
rect 1562 530 1596 706
rect 1720 530 1754 706
rect -1266 324 -1232 400
rect -1108 324 -1074 400
rect 1636 406 1672 440
rect -1346 174 -1308 210
rect -1188 172 -1150 206
rect 498 164 532 340
rect 656 164 690 340
rect 814 164 848 340
rect 1562 154 1596 330
rect 1720 154 1754 330
rect 574 80 610 114
rect 730 80 766 114
rect -2460 -628 -1922 -231
rect -1642 -520 -1608 -444
rect -1484 -520 -1450 -444
rect -1326 -520 -1292 -444
rect -1428 -622 -1388 -582
rect -2602 -858 -2558 -774
rect -2460 -1389 -1922 -992
rect -1196 -1324 -1162 -448
rect -1038 -1324 -1004 -448
rect -880 -1324 -846 -448
rect -1328 -1414 -1288 -1374
rect -1174 -1420 -1128 -1386
rect -2460 -1924 -1922 -1527
rect -1266 -2042 -1232 -1866
rect -1108 -2042 -1074 -1866
rect -978 -2042 -944 -1982
rect -820 -2042 -786 -1982
rect -2388 -2204 -2344 -2120
rect -1048 -2160 -1010 -2124
rect -1424 -2630 -1390 -2554
rect -1266 -2630 -1232 -2554
rect -1108 -2630 -1074 -2554
rect -1348 -2782 -1310 -2746
rect -1190 -2784 -1152 -2748
<< metal1 >>
rect -1304 5558 -1240 5564
rect -1304 5544 -1298 5558
rect -1490 5506 -1298 5544
rect -1246 5544 -1240 5558
rect -1246 5506 -840 5544
rect -1490 5504 -840 5506
rect -1648 5460 -1602 5472
rect -1648 5384 -1642 5460
rect -1608 5384 -1602 5460
rect -1648 5372 -1602 5384
rect -1490 5460 -1444 5504
rect -1304 5500 -1240 5504
rect -1490 5384 -1484 5460
rect -1450 5384 -1444 5460
rect -1490 5372 -1444 5384
rect -1332 5460 -1286 5472
rect -1332 5384 -1326 5460
rect -1292 5384 -1286 5460
rect -1440 5328 -1376 5334
rect -1440 5276 -1434 5328
rect -1382 5276 -1376 5328
rect -1440 5270 -1376 5276
rect -1332 4542 -1286 5384
rect -1202 5456 -1156 5504
rect -1202 4580 -1196 5456
rect -1162 4580 -1156 5456
rect -1202 4568 -1156 4580
rect -1044 5456 -998 5468
rect -1044 4580 -1038 5456
rect -1004 4580 -998 5456
rect -1340 4536 -1276 4542
rect -1340 4484 -1334 4536
rect -1282 4524 -1276 4536
rect -1282 4518 -1116 4524
rect -1282 4484 -1174 4518
rect -1128 4484 -1116 4518
rect -1340 4478 -1116 4484
rect -1044 4128 -998 4580
rect -886 5456 -840 5504
rect -886 4580 -880 5456
rect -846 4580 -840 5456
rect -886 4568 -840 4580
rect -784 4128 -720 4134
rect -1044 4078 -778 4128
rect -826 4076 -778 4078
rect -726 4076 -720 4128
rect -826 4070 -720 4076
rect -1272 4038 -1226 4050
rect -1272 3862 -1266 4038
rect -1232 3862 -1226 4038
rect -2270 3238 -2108 3842
rect -1858 3796 -1794 3802
rect -1858 3744 -1852 3796
rect -1800 3744 -1794 3796
rect -1858 3738 -1794 3744
rect -1444 3350 -1376 3362
rect -1444 3284 -1434 3350
rect -1382 3284 -1376 3350
rect -1272 3350 -1226 3862
rect -1114 4038 -1068 4050
rect -1114 3862 -1108 4038
rect -1074 3894 -1068 4038
rect -984 3922 -938 3934
rect -984 3894 -978 3922
rect -1074 3882 -978 3894
rect -1074 3862 -1052 3882
rect -1114 3850 -1052 3862
rect -1058 3830 -1052 3850
rect -1000 3862 -978 3882
rect -944 3862 -938 3922
rect -1000 3850 -938 3862
rect -826 3922 -780 4070
rect -826 3862 -820 3922
rect -786 3862 -780 3922
rect -826 3850 -780 3862
rect -1000 3830 -994 3850
rect -1058 3824 -994 3830
rect -894 3812 -714 3814
rect -894 3806 -708 3812
rect -894 3802 -766 3806
rect -894 3766 -882 3802
rect -844 3766 -766 3802
rect -894 3754 -766 3766
rect -714 3754 -708 3806
rect -894 3748 -708 3754
rect -1430 3274 -1424 3284
rect -1390 3274 -1384 3284
rect -1430 3262 -1384 3274
rect -1272 3274 -1266 3350
rect -1232 3274 -1226 3350
rect -1126 3350 -1058 3362
rect -1126 3342 -1108 3350
rect -1074 3342 -1058 3350
rect -1126 3290 -1116 3342
rect -1064 3290 -1058 3342
rect -1126 3284 -1108 3290
rect -1272 3262 -1226 3274
rect -1114 3274 -1108 3284
rect -1074 3284 -1058 3290
rect -1074 3274 -1068 3284
rect -1114 3262 -1068 3274
rect -2470 3232 -1908 3238
rect -2470 2835 -2458 3232
rect -1920 2835 -1908 3232
rect -1462 3166 -1296 3172
rect -1462 3114 -1456 3166
rect -1404 3160 -1296 3166
rect -1404 3124 -1346 3160
rect -1308 3124 -1296 3160
rect -1404 3114 -1296 3124
rect -1462 3108 -1296 3114
rect -1202 3156 -1140 3168
rect -1202 3120 -1190 3156
rect -1152 3120 -1140 3156
rect -1202 3012 -1140 3120
rect -2470 2829 -1908 2835
rect -1782 2952 -1140 3012
rect -2470 2697 -1908 2703
rect -2470 2300 -2458 2697
rect -1920 2300 -1908 2697
rect -2470 2294 -1908 2300
rect -2626 2160 -2534 2226
rect -2626 2076 -2602 2160
rect -2558 2076 -2534 2160
rect -2626 694 -2534 2076
rect -2268 2152 -2110 2294
rect -1782 2152 -1722 2952
rect 1628 2678 1694 2684
rect 1628 2632 1634 2678
rect 1480 2626 1634 2632
rect 1688 2632 1694 2678
rect 2528 2678 2594 2684
rect 2528 2632 2534 2678
rect 1688 2626 1842 2632
rect -1304 2612 -1240 2618
rect -1304 2594 -1298 2612
rect -1490 2560 -1298 2594
rect -1246 2594 -1240 2612
rect -1246 2560 -840 2594
rect -1490 2554 -840 2560
rect -1648 2510 -1602 2522
rect -1648 2434 -1642 2510
rect -1608 2434 -1602 2510
rect -1648 2422 -1602 2434
rect -1490 2510 -1444 2554
rect -1490 2434 -1484 2510
rect -1450 2434 -1444 2510
rect -1490 2422 -1444 2434
rect -1332 2510 -1286 2522
rect -1332 2434 -1326 2510
rect -1292 2434 -1286 2510
rect -1440 2378 -1376 2384
rect -1440 2326 -1434 2378
rect -1382 2326 -1376 2378
rect -1440 2320 -1376 2326
rect -2268 2092 -1720 2152
rect -2268 1950 -2110 2092
rect -2470 1944 -1908 1950
rect -2470 1547 -2458 1944
rect -1920 1547 -1908 1944
rect -1332 1592 -1286 2434
rect -1202 2506 -1156 2554
rect -1202 1630 -1196 2506
rect -1162 1630 -1156 2506
rect -1202 1618 -1156 1630
rect -1044 2506 -998 2518
rect -1044 1630 -1038 2506
rect -1004 1630 -998 2506
rect -2470 1541 -1908 1547
rect -1340 1586 -1276 1592
rect -1340 1534 -1334 1586
rect -1282 1574 -1276 1586
rect -1282 1568 -1116 1574
rect -1282 1534 -1174 1568
rect -1128 1534 -1116 1568
rect -1340 1528 -1116 1534
rect -2470 1265 -1908 1271
rect -2470 868 -2458 1265
rect -1920 868 -1908 1265
rect -1044 1178 -998 1630
rect -886 2506 -840 2554
rect -886 1630 -880 2506
rect -846 1630 -840 2506
rect 1480 2592 1842 2626
rect 1480 2538 1526 2592
rect 1480 2362 1486 2538
rect 1520 2362 1526 2538
rect 1480 2350 1526 2362
rect 1638 2538 1684 2550
rect 1638 2362 1644 2538
rect 1678 2362 1684 2538
rect 1638 2308 1684 2362
rect 1796 2538 1842 2592
rect 1796 2362 1802 2538
rect 1836 2362 1842 2538
rect 1796 2350 1842 2362
rect 2380 2626 2534 2632
rect 2588 2632 2594 2678
rect 2588 2626 2742 2632
rect 2380 2592 2742 2626
rect 2380 2538 2426 2592
rect 2380 2362 2386 2538
rect 2420 2362 2426 2538
rect 2380 2350 2426 2362
rect 2538 2538 2584 2550
rect 2538 2362 2544 2538
rect 2578 2362 2584 2538
rect 1858 2312 1922 2318
rect 1858 2308 1864 2312
rect 1480 2264 1864 2308
rect 1480 2204 1526 2264
rect 1858 2260 1864 2264
rect 1916 2260 1922 2312
rect 2538 2308 2584 2362
rect 2696 2538 2742 2592
rect 2696 2362 2702 2538
rect 2736 2362 2742 2538
rect 3442 2570 3488 2582
rect 3442 2420 3448 2570
rect 2696 2350 2742 2362
rect 3432 2414 3448 2420
rect 3482 2420 3488 2570
rect 3600 2570 3646 2582
rect 3482 2414 3498 2420
rect 3432 2362 3438 2414
rect 3492 2362 3498 2414
rect 3432 2356 3498 2362
rect 3600 2394 3606 2570
rect 3640 2394 3646 2570
rect 3442 2338 3488 2356
rect 3600 2350 3646 2394
rect 3600 2344 3702 2350
rect 2758 2312 2822 2318
rect 2758 2308 2764 2312
rect 1858 2254 1922 2260
rect 2380 2264 2764 2308
rect 640 2162 706 2168
rect 640 2116 646 2162
rect 492 2110 646 2116
rect 700 2116 706 2162
rect 700 2110 854 2116
rect 492 2076 854 2110
rect 492 2022 538 2076
rect 492 1846 498 2022
rect 532 1846 538 2022
rect 492 1834 538 1846
rect 650 2022 696 2034
rect 650 1846 656 2022
rect 690 1846 696 2022
rect 650 1792 696 1846
rect 808 2022 854 2076
rect 808 1846 814 2022
rect 848 1846 854 2022
rect 1480 2028 1486 2204
rect 1520 2028 1526 2204
rect 1480 2016 1526 2028
rect 1638 2204 1684 2216
rect 1638 2028 1644 2204
rect 1678 2028 1684 2204
rect 1638 2016 1684 2028
rect 1796 2204 1842 2216
rect 1796 2028 1802 2204
rect 1836 2028 1842 2204
rect 1796 2024 1842 2028
rect 2380 2204 2426 2264
rect 2758 2260 2764 2264
rect 2816 2260 2822 2312
rect 2758 2254 2822 2260
rect 3508 2312 3572 2318
rect 3508 2260 3514 2312
rect 3566 2260 3572 2312
rect 3508 2254 3572 2260
rect 3600 2292 3644 2344
rect 3696 2292 3702 2344
rect 3600 2286 3702 2292
rect 2380 2028 2386 2204
rect 2420 2028 2426 2204
rect 1796 2018 1868 2024
rect 1548 1986 1612 1992
rect 1548 1934 1554 1986
rect 1606 1934 1612 1986
rect 1548 1928 1612 1934
rect 1704 1986 1768 1992
rect 1704 1934 1710 1986
rect 1762 1934 1768 1986
rect 1796 1966 1808 2018
rect 1862 1966 1868 2018
rect 2380 2016 2426 2028
rect 2538 2204 2584 2216
rect 2538 2028 2544 2204
rect 2578 2028 2584 2204
rect 2538 2016 2584 2028
rect 2696 2204 2742 2216
rect 2696 2028 2702 2204
rect 2736 2036 2742 2204
rect 3442 2194 3488 2206
rect 2736 2030 2768 2036
rect 1796 1960 1868 1966
rect 2448 1986 2512 1992
rect 1704 1928 1768 1934
rect 2448 1934 2454 1986
rect 2506 1934 2512 1986
rect 2448 1928 2512 1934
rect 2604 1986 2668 1992
rect 2604 1934 2610 1986
rect 2662 1934 2668 1986
rect 2696 1978 2708 2028
rect 2762 1978 2768 2030
rect 3442 2018 3448 2194
rect 3482 2018 3488 2194
rect 2696 1972 2768 1978
rect 3300 2012 3366 2014
rect 3442 2012 3488 2018
rect 3600 2194 3646 2286
rect 3600 2018 3606 2194
rect 3640 2018 3646 2194
rect 3300 2008 3498 2012
rect 3300 1956 3306 2008
rect 3360 1956 3498 2008
rect 3600 2006 3646 2018
rect 3300 1952 3498 1956
rect 3300 1950 3366 1952
rect 2604 1928 2668 1934
rect 808 1834 854 1846
rect 870 1796 934 1802
rect 870 1792 876 1796
rect -886 1618 -840 1630
rect 492 1748 876 1792
rect 492 1688 538 1748
rect 870 1744 876 1748
rect 928 1744 934 1796
rect 870 1738 934 1744
rect 1628 1776 1694 1782
rect 1628 1730 1634 1776
rect 1480 1724 1634 1730
rect 1688 1730 1694 1776
rect 1688 1724 1842 1730
rect 492 1512 498 1688
rect 532 1512 538 1688
rect 492 1500 538 1512
rect 650 1688 696 1700
rect 650 1512 656 1688
rect 690 1512 696 1688
rect 650 1500 696 1512
rect 808 1688 854 1700
rect 808 1512 814 1688
rect 848 1514 854 1688
rect 1480 1690 1842 1724
rect 1480 1636 1526 1690
rect 848 1512 880 1514
rect 808 1508 880 1512
rect 562 1470 626 1476
rect 6 1456 72 1462
rect 6 1404 12 1456
rect 66 1404 72 1456
rect 562 1418 568 1470
rect 620 1418 626 1470
rect 562 1412 626 1418
rect 716 1470 780 1476
rect 716 1418 722 1470
rect 774 1418 780 1470
rect 808 1456 820 1508
rect 874 1456 880 1508
rect 814 1450 880 1456
rect 1480 1460 1486 1636
rect 1520 1460 1526 1636
rect 1480 1448 1526 1460
rect 1638 1636 1684 1648
rect 1638 1460 1644 1636
rect 1678 1460 1684 1636
rect 716 1412 780 1418
rect 1638 1406 1684 1460
rect 1796 1636 1842 1690
rect 1796 1460 1802 1636
rect 1836 1460 1842 1636
rect 2528 1620 2594 1626
rect 2528 1574 2534 1620
rect 1796 1448 1842 1460
rect 2376 1568 2534 1574
rect 2588 1574 2594 1620
rect 2588 1568 2738 1574
rect 2376 1534 2738 1568
rect 2376 1480 2422 1534
rect 1858 1410 1922 1416
rect 1858 1406 1864 1410
rect 6 1396 72 1404
rect 1480 1362 1864 1406
rect 1480 1302 1526 1362
rect 1858 1358 1864 1362
rect 1916 1358 1922 1410
rect 1858 1352 1922 1358
rect -784 1178 -720 1184
rect -1044 1128 -778 1178
rect -826 1126 -778 1128
rect -726 1126 -720 1178
rect -826 1120 -720 1126
rect 1480 1126 1486 1302
rect 1520 1126 1526 1302
rect -2470 862 -1908 868
rect -1272 1088 -1226 1100
rect -1272 912 -1266 1088
rect -1232 912 -1226 1088
rect -2626 610 -2602 694
rect -2558 610 -2534 694
rect -2626 -774 -2534 610
rect -2270 680 -2108 862
rect -2270 620 -1720 680
rect -2270 454 -2108 620
rect -2472 448 -1910 454
rect -2472 51 -2460 448
rect -1922 51 -1910 448
rect -2472 45 -1910 51
rect -1782 72 -1720 620
rect -1444 400 -1376 412
rect -1444 334 -1434 400
rect -1382 334 -1376 400
rect -1272 400 -1226 912
rect -1114 1088 -1068 1100
rect -1114 912 -1108 1088
rect -1074 944 -1068 1088
rect -984 972 -938 984
rect -984 944 -978 972
rect -1074 932 -978 944
rect -1074 912 -1052 932
rect -1114 900 -1052 912
rect -1058 880 -1052 900
rect -1000 912 -978 932
rect -944 912 -938 972
rect -1000 900 -938 912
rect -826 972 -780 1120
rect 1480 1114 1526 1126
rect 1638 1302 1684 1314
rect 1638 1126 1644 1302
rect 1678 1126 1684 1302
rect 1638 1114 1684 1126
rect 1796 1302 1842 1314
rect 1796 1126 1802 1302
rect 1836 1126 1842 1302
rect 2376 1304 2382 1480
rect 2416 1304 2422 1480
rect 2376 1292 2422 1304
rect 2534 1480 2580 1492
rect 2534 1304 2540 1480
rect 2574 1304 2580 1480
rect 2534 1250 2580 1304
rect 2692 1480 2738 1534
rect 2692 1304 2698 1480
rect 2732 1304 2738 1480
rect 3442 1512 3488 1524
rect 3442 1360 3448 1512
rect 2692 1292 2738 1304
rect 3432 1354 3448 1360
rect 3482 1360 3488 1512
rect 3600 1512 3646 1524
rect 3482 1354 3498 1360
rect 3432 1302 3438 1354
rect 3492 1302 3498 1354
rect 3432 1296 3498 1302
rect 3600 1336 3606 1512
rect 3640 1336 3646 1512
rect 3442 1280 3488 1296
rect 3600 1288 3646 1336
rect 3600 1282 3702 1288
rect 2754 1254 2818 1260
rect 2754 1250 2760 1254
rect 1796 1122 1842 1126
rect 2376 1206 2760 1250
rect 2376 1146 2422 1206
rect 2754 1202 2760 1206
rect 2812 1202 2818 1254
rect 2754 1196 2818 1202
rect 3508 1254 3572 1260
rect 3508 1202 3514 1254
rect 3566 1202 3572 1254
rect 3508 1196 3572 1202
rect 3600 1230 3644 1282
rect 3696 1230 3702 1282
rect 3600 1224 3702 1230
rect 1796 1116 1868 1122
rect 1548 1084 1612 1090
rect 1548 1032 1554 1084
rect 1606 1032 1612 1084
rect 1548 1026 1612 1032
rect 1704 1084 1768 1090
rect 1704 1032 1710 1084
rect 1762 1032 1768 1084
rect 1796 1070 1808 1116
rect 1802 1064 1808 1070
rect 1862 1064 1868 1116
rect 1802 1058 1868 1064
rect 1704 1026 1768 1032
rect -826 912 -820 972
rect -786 912 -780 972
rect 2376 970 2382 1146
rect 2416 970 2422 1146
rect 2376 958 2422 970
rect 2534 1146 2580 1158
rect 2534 970 2540 1146
rect 2574 970 2580 1146
rect 2534 958 2580 970
rect 2692 1146 2738 1158
rect 2692 970 2698 1146
rect 2732 972 2738 1146
rect 3442 1136 3488 1148
rect 2732 970 2764 972
rect 2692 966 2764 970
rect -826 900 -780 912
rect 2444 928 2508 934
rect -1000 880 -994 900
rect -1058 874 -994 880
rect 2444 876 2450 928
rect 2502 876 2508 928
rect 6 866 72 872
rect 2444 870 2508 876
rect 2600 928 2664 934
rect 2600 876 2606 928
rect 2658 876 2664 928
rect 2692 914 2704 966
rect 2758 914 2764 966
rect 3442 960 3448 1136
rect 3482 960 3488 1136
rect 3442 954 3488 960
rect 3600 1136 3646 1224
rect 3600 960 3606 1136
rect 3640 960 3646 1136
rect 3438 952 3498 954
rect 2698 908 2764 914
rect 3432 946 3498 952
rect 3600 948 3646 960
rect 3432 894 3438 946
rect 3492 894 3498 946
rect 3432 888 3498 894
rect 2600 870 2664 876
rect -912 854 -850 866
rect -912 818 -900 854
rect -862 818 -850 854
rect -912 716 -850 818
rect 6 814 12 866
rect 66 814 72 866
rect 6 806 72 814
rect 640 814 706 820
rect 640 768 646 814
rect 492 762 646 768
rect 700 768 706 814
rect 700 762 854 768
rect 492 728 854 762
rect -772 716 -708 722
rect -912 664 -766 716
rect -714 664 -708 716
rect -772 658 -708 664
rect 492 674 538 728
rect 492 498 498 674
rect 532 498 538 674
rect 492 486 538 498
rect 650 674 696 686
rect 650 498 656 674
rect 690 498 696 674
rect 650 444 696 498
rect 808 674 854 728
rect 808 498 814 674
rect 848 498 854 674
rect 1556 706 1602 718
rect 1556 554 1562 706
rect 808 486 854 498
rect 1544 548 1562 554
rect 1596 554 1602 706
rect 1714 706 1760 718
rect 1596 548 1610 554
rect 1544 496 1550 548
rect 1604 496 1610 548
rect 1544 490 1610 496
rect 1714 530 1720 706
rect 1754 530 1760 706
rect 1556 474 1602 490
rect 1714 486 1760 530
rect 1714 480 1820 486
rect 870 448 934 454
rect 870 444 876 448
rect -1430 324 -1424 334
rect -1390 324 -1384 334
rect -1430 312 -1384 324
rect -1272 324 -1266 400
rect -1232 324 -1226 400
rect -1126 400 -1058 412
rect -1126 392 -1108 400
rect -1074 392 -1058 400
rect -1126 340 -1116 392
rect -1064 340 -1058 392
rect -1126 334 -1108 340
rect -1272 312 -1226 324
rect -1114 324 -1108 334
rect -1074 334 -1058 340
rect 492 400 876 444
rect 492 340 538 400
rect 870 396 876 400
rect 928 396 934 448
rect 870 390 934 396
rect 1622 448 1686 454
rect 1622 396 1628 448
rect 1680 396 1686 448
rect 1622 390 1686 396
rect 1714 428 1762 480
rect 1814 428 1820 480
rect 1714 422 1820 428
rect -1074 324 -1068 334
rect -1114 312 -1068 324
rect -1462 216 -1296 222
rect -1462 164 -1456 216
rect -1404 210 -1296 216
rect -1404 174 -1346 210
rect -1308 174 -1296 210
rect -1404 164 -1296 174
rect -1462 158 -1296 164
rect -1200 206 -1138 224
rect -1200 172 -1188 206
rect -1150 172 -1138 206
rect -1200 72 -1138 172
rect 492 164 498 340
rect 532 164 538 340
rect 492 152 538 164
rect 650 340 696 352
rect 650 164 656 340
rect 690 164 696 340
rect 650 152 696 164
rect 808 340 854 352
rect 808 164 814 340
rect 848 164 854 340
rect 808 162 854 164
rect 1556 330 1602 342
rect 808 156 880 162
rect -1782 12 -1138 72
rect 560 122 624 128
rect 560 70 566 122
rect 618 70 624 122
rect 560 64 624 70
rect 716 122 780 128
rect 716 70 722 122
rect 774 70 780 122
rect 808 108 820 156
rect 814 104 820 108
rect 874 104 880 156
rect 1556 154 1562 330
rect 1596 154 1602 330
rect 1556 148 1602 154
rect 1714 330 1760 422
rect 1714 154 1720 330
rect 1754 154 1760 330
rect 814 98 880 104
rect 1546 142 1612 148
rect 1714 142 1760 154
rect 1546 90 1552 142
rect 1606 90 1612 142
rect 1546 84 1612 90
rect 716 64 780 70
rect -2472 -231 -1910 -225
rect -2472 -628 -2460 -231
rect -1922 -628 -1910 -231
rect -1304 -346 -1240 -340
rect -1304 -360 -1298 -346
rect -1490 -398 -1298 -360
rect -1246 -360 -1240 -346
rect -1246 -398 -840 -360
rect -1490 -400 -840 -398
rect -1648 -444 -1602 -432
rect -1648 -520 -1642 -444
rect -1608 -520 -1602 -444
rect -1648 -532 -1602 -520
rect -1490 -444 -1444 -400
rect -1304 -404 -1240 -400
rect -1490 -520 -1484 -444
rect -1450 -520 -1444 -444
rect -1490 -532 -1444 -520
rect -1332 -444 -1286 -432
rect -1332 -520 -1326 -444
rect -1292 -520 -1286 -444
rect -2472 -634 -1910 -628
rect -1440 -576 -1376 -570
rect -1440 -628 -1434 -576
rect -1382 -628 -1376 -576
rect -1440 -634 -1376 -628
rect -2626 -858 -2602 -774
rect -2558 -858 -2534 -774
rect -2626 -2096 -2534 -858
rect -2270 -786 -2108 -634
rect -2270 -846 -1720 -786
rect -2270 -986 -2108 -846
rect -2472 -992 -1910 -986
rect -2472 -1389 -2460 -992
rect -1922 -1389 -1910 -992
rect -2472 -1395 -1910 -1389
rect -2472 -1527 -1910 -1521
rect -2472 -1924 -2460 -1527
rect -1922 -1924 -1910 -1527
rect -2472 -1930 -1910 -1924
rect -2626 -2114 -2320 -2096
rect -2270 -2114 -2108 -1930
rect -2626 -2120 -2108 -2114
rect -2626 -2204 -2388 -2120
rect -2344 -2204 -2108 -2120
rect -2626 -2210 -2108 -2204
rect -2626 -2228 -2320 -2210
rect -2270 -2286 -2108 -2210
rect -2270 -2410 -2242 -2286
rect -2132 -2410 -2108 -2286
rect -2270 -2432 -2108 -2410
rect -1782 -2868 -1720 -846
rect -1332 -1362 -1286 -520
rect -1202 -448 -1156 -400
rect -1202 -1324 -1196 -448
rect -1162 -1324 -1156 -448
rect -1202 -1336 -1156 -1324
rect -1044 -448 -998 -436
rect -1044 -1324 -1038 -448
rect -1004 -1324 -998 -448
rect -1340 -1368 -1276 -1362
rect -1340 -1420 -1334 -1368
rect -1282 -1380 -1276 -1368
rect -1282 -1386 -1116 -1380
rect -1282 -1420 -1174 -1386
rect -1128 -1420 -1116 -1386
rect -1340 -1426 -1116 -1420
rect -1044 -1776 -998 -1324
rect -886 -448 -840 -400
rect -886 -1324 -880 -448
rect -846 -1324 -840 -448
rect -886 -1336 -840 -1324
rect -784 -1776 -720 -1770
rect -1044 -1826 -778 -1776
rect -826 -1828 -778 -1826
rect -726 -1828 -720 -1776
rect -826 -1834 -720 -1828
rect -1272 -1866 -1226 -1854
rect -1272 -2042 -1266 -1866
rect -1232 -2042 -1226 -1866
rect -1444 -2554 -1376 -2542
rect -1444 -2620 -1434 -2554
rect -1382 -2620 -1376 -2554
rect -1272 -2554 -1226 -2042
rect -1114 -1866 -1068 -1854
rect -1114 -2042 -1108 -1866
rect -1074 -2010 -1068 -1866
rect -984 -1982 -938 -1970
rect -984 -2010 -978 -1982
rect -1074 -2022 -978 -2010
rect -1074 -2042 -1052 -2022
rect -1114 -2054 -1052 -2042
rect -1058 -2074 -1052 -2054
rect -1000 -2042 -978 -2022
rect -944 -2042 -938 -1982
rect -1000 -2054 -938 -2042
rect -826 -1982 -780 -1834
rect -826 -2042 -820 -1982
rect -786 -2042 -780 -1982
rect -826 -2054 -780 -2042
rect -1000 -2074 -994 -2054
rect -1058 -2080 -994 -2074
rect -1060 -2124 -998 -2112
rect -1060 -2160 -1048 -2124
rect -1010 -2160 -998 -2124
rect -1060 -2164 -998 -2160
rect -1062 -2170 -998 -2164
rect -1062 -2222 -1056 -2170
rect -1004 -2222 -998 -2170
rect -1062 -2228 -998 -2222
rect -772 -2358 -708 -2352
rect -772 -2410 -766 -2358
rect -714 -2410 -708 -2358
rect -772 -2416 -708 -2410
rect -1430 -2630 -1424 -2620
rect -1390 -2630 -1384 -2620
rect -1430 -2642 -1384 -2630
rect -1272 -2630 -1266 -2554
rect -1232 -2630 -1226 -2554
rect -1126 -2554 -1058 -2542
rect -1126 -2562 -1108 -2554
rect -1074 -2562 -1058 -2554
rect -1126 -2614 -1116 -2562
rect -1064 -2614 -1058 -2562
rect -1126 -2620 -1108 -2614
rect -1272 -2642 -1226 -2630
rect -1114 -2630 -1108 -2620
rect -1074 -2620 -1058 -2614
rect -1074 -2630 -1068 -2620
rect -1114 -2642 -1068 -2630
rect -1360 -2738 -1296 -2732
rect -1360 -2790 -1354 -2738
rect -1302 -2790 -1296 -2738
rect -1360 -2796 -1296 -2790
rect -1202 -2748 -1140 -2736
rect -1202 -2784 -1190 -2748
rect -1152 -2784 -1140 -2748
rect -1360 -2800 -1298 -2796
rect -1202 -2868 -1140 -2784
rect -1782 -2928 -1140 -2868
<< via1 >>
rect -1298 5506 -1246 5558
rect -1434 5322 -1382 5328
rect -1434 5282 -1428 5322
rect -1428 5282 -1388 5322
rect -1388 5282 -1382 5322
rect -1434 5276 -1382 5282
rect -1334 4530 -1282 4536
rect -1334 4490 -1328 4530
rect -1328 4490 -1288 4530
rect -1288 4490 -1282 4530
rect -1334 4484 -1282 4490
rect -778 4076 -726 4128
rect -1852 3744 -1800 3796
rect -1434 3284 -1424 3350
rect -1424 3284 -1390 3350
rect -1390 3284 -1382 3350
rect -1052 3830 -1000 3882
rect -766 3754 -714 3806
rect -1116 3290 -1108 3342
rect -1108 3290 -1074 3342
rect -1074 3290 -1064 3342
rect -1456 3114 -1404 3166
rect 1634 2626 1688 2678
rect -1298 2560 -1246 2612
rect -1434 2372 -1382 2378
rect -1434 2332 -1428 2372
rect -1428 2332 -1388 2372
rect -1388 2332 -1382 2372
rect -1434 2326 -1382 2332
rect -1334 1580 -1282 1586
rect -1334 1540 -1328 1580
rect -1328 1540 -1288 1580
rect -1288 1540 -1282 1580
rect -1334 1534 -1282 1540
rect 2534 2626 2588 2678
rect 1864 2260 1916 2312
rect 3438 2394 3448 2414
rect 3448 2394 3482 2414
rect 3482 2394 3492 2414
rect 3438 2362 3492 2394
rect 646 2110 700 2162
rect 2764 2260 2816 2312
rect 3514 2304 3566 2312
rect 3514 2270 3522 2304
rect 3522 2270 3558 2304
rect 3558 2270 3566 2304
rect 3514 2260 3566 2270
rect 3644 2292 3696 2344
rect 1554 1978 1606 1986
rect 1554 1944 1562 1978
rect 1562 1944 1598 1978
rect 1598 1944 1606 1978
rect 1554 1934 1606 1944
rect 1710 1978 1762 1986
rect 1710 1944 1718 1978
rect 1718 1944 1754 1978
rect 1754 1944 1762 1978
rect 1710 1934 1762 1944
rect 1808 1966 1862 2018
rect 2708 2028 2736 2030
rect 2736 2028 2762 2030
rect 2454 1978 2506 1986
rect 2454 1944 2462 1978
rect 2462 1944 2498 1978
rect 2498 1944 2506 1978
rect 2454 1934 2506 1944
rect 2610 1978 2662 1986
rect 2610 1944 2618 1978
rect 2618 1944 2654 1978
rect 2654 1944 2662 1978
rect 2610 1934 2662 1944
rect 2708 1978 2762 2028
rect 3306 1956 3360 2008
rect 876 1744 928 1796
rect 1634 1724 1688 1776
rect 12 1404 66 1456
rect 568 1462 620 1470
rect 568 1428 576 1462
rect 576 1428 612 1462
rect 612 1428 620 1462
rect 568 1418 620 1428
rect 722 1462 774 1470
rect 722 1428 730 1462
rect 730 1428 766 1462
rect 766 1428 774 1462
rect 722 1418 774 1428
rect 820 1456 874 1508
rect 2534 1568 2588 1620
rect 1864 1358 1916 1410
rect -778 1126 -726 1178
rect -1434 334 -1424 400
rect -1424 334 -1390 400
rect -1390 334 -1382 400
rect -1052 880 -1000 932
rect 3438 1336 3448 1354
rect 3448 1336 3482 1354
rect 3482 1336 3492 1354
rect 3438 1302 3492 1336
rect 2760 1202 2812 1254
rect 3514 1246 3566 1254
rect 3514 1212 3522 1246
rect 3522 1212 3558 1246
rect 3558 1212 3566 1246
rect 3514 1202 3566 1212
rect 3644 1230 3696 1282
rect 1554 1076 1606 1084
rect 1554 1042 1562 1076
rect 1562 1042 1598 1076
rect 1598 1042 1606 1076
rect 1554 1032 1606 1042
rect 1710 1076 1762 1084
rect 1710 1042 1718 1076
rect 1718 1042 1754 1076
rect 1754 1042 1762 1076
rect 1710 1032 1762 1042
rect 1808 1064 1862 1116
rect 2450 920 2502 928
rect 2450 886 2458 920
rect 2458 886 2494 920
rect 2494 886 2502 920
rect 2450 876 2502 886
rect 2606 920 2658 928
rect 2606 886 2614 920
rect 2614 886 2650 920
rect 2650 886 2658 920
rect 2606 876 2658 886
rect 2704 914 2758 966
rect 3438 894 3492 946
rect 12 814 66 866
rect 646 762 700 814
rect -766 664 -714 716
rect 1550 530 1562 548
rect 1562 530 1596 548
rect 1596 530 1604 548
rect 1550 496 1604 530
rect -1116 340 -1108 392
rect -1108 340 -1074 392
rect -1074 340 -1064 392
rect 876 396 928 448
rect 1628 440 1680 448
rect 1628 406 1636 440
rect 1636 406 1672 440
rect 1672 406 1680 440
rect 1628 396 1680 406
rect 1762 428 1814 480
rect -1456 164 -1404 216
rect 566 114 618 122
rect 566 80 574 114
rect 574 80 610 114
rect 610 80 618 114
rect 566 70 618 80
rect 722 114 774 122
rect 722 80 730 114
rect 730 80 766 114
rect 766 80 774 114
rect 722 70 774 80
rect 820 104 874 156
rect 1552 90 1606 142
rect -1298 -398 -1246 -346
rect -1434 -582 -1382 -576
rect -1434 -622 -1428 -582
rect -1428 -622 -1388 -582
rect -1388 -622 -1382 -582
rect -1434 -628 -1382 -622
rect -2242 -2410 -2132 -2286
rect -1334 -1374 -1282 -1368
rect -1334 -1414 -1328 -1374
rect -1328 -1414 -1288 -1374
rect -1288 -1414 -1282 -1374
rect -1334 -1420 -1282 -1414
rect -778 -1828 -726 -1776
rect -1434 -2620 -1424 -2554
rect -1424 -2620 -1390 -2554
rect -1390 -2620 -1382 -2554
rect -1052 -2074 -1000 -2022
rect -1056 -2222 -1004 -2170
rect -766 -2410 -714 -2358
rect -1116 -2614 -1108 -2562
rect -1108 -2614 -1074 -2562
rect -1074 -2614 -1064 -2562
rect -1354 -2746 -1302 -2738
rect -1354 -2782 -1348 -2746
rect -1348 -2782 -1310 -2746
rect -1310 -2782 -1302 -2746
rect -1354 -2790 -1302 -2782
<< metal2 >>
rect -1310 5560 -1234 5570
rect -1310 5504 -1300 5560
rect -1244 5504 -1234 5560
rect -1310 5494 -1234 5504
rect -1440 5328 -1376 5334
rect -1440 5276 -1434 5328
rect -1382 5276 -1376 5328
rect -1440 5270 -1376 5276
rect -1864 3798 -1788 3808
rect -1864 3742 -1854 3798
rect -1798 3742 -1788 3798
rect -1864 3732 -1788 3742
rect -1436 3362 -1380 5270
rect -1340 4536 -1276 4542
rect -1340 4484 -1334 4536
rect -1282 4484 -1276 4536
rect -1340 4478 -1276 4484
rect -1334 3456 -1282 4478
rect -784 4128 -720 4134
rect -784 4076 -778 4128
rect -726 4126 -720 4128
rect -726 4078 -162 4126
rect -726 4076 -720 4078
rect -784 4070 -720 4076
rect -1064 3884 -988 3894
rect -1064 3828 -1054 3884
rect -998 3828 -988 3884
rect -1064 3818 -988 3828
rect -778 3808 -702 3818
rect -778 3752 -768 3808
rect -712 3752 -702 3808
rect -778 3742 -702 3752
rect -1334 3404 -1064 3456
rect -1116 3362 -1064 3404
rect -1444 3350 -1376 3362
rect -1444 3284 -1434 3350
rect -1382 3284 -1376 3350
rect -1126 3342 -1058 3362
rect -1126 3290 -1116 3342
rect -1064 3290 -1058 3342
rect -1126 3284 -1058 3290
rect -1468 3168 -1392 3178
rect -1468 3112 -1458 3168
rect -1402 3112 -1392 3168
rect -1468 3102 -1392 3112
rect -1310 2614 -1234 2624
rect -1310 2558 -1300 2614
rect -1244 2558 -1234 2614
rect -1310 2548 -1234 2558
rect -1440 2378 -1376 2384
rect -1440 2326 -1434 2378
rect -1382 2326 -1376 2378
rect -1440 2320 -1376 2326
rect -1436 412 -1380 2320
rect -1340 1586 -1276 1592
rect -1340 1534 -1334 1586
rect -1282 1534 -1276 1586
rect -1340 1528 -1276 1534
rect -1334 506 -1282 1528
rect -210 1326 -162 4078
rect 1622 2680 1700 2690
rect 1622 2624 1632 2680
rect 1690 2624 1700 2680
rect 1622 2612 1700 2624
rect 2522 2680 2600 2690
rect 2522 2624 2532 2680
rect 2590 2624 2600 2680
rect 2522 2612 2600 2624
rect 3426 2416 3504 2426
rect 3426 2360 3436 2416
rect 3494 2360 3504 2416
rect 3426 2348 3504 2360
rect 3638 2344 3702 2350
rect 1858 2312 1922 2318
rect 1858 2260 1864 2312
rect 1916 2306 1922 2312
rect 2758 2312 2822 2318
rect 1916 2266 2348 2306
rect 1916 2260 1922 2266
rect 1858 2254 1922 2260
rect 634 2164 712 2174
rect 634 2108 644 2164
rect 702 2108 712 2164
rect 634 2096 712 2108
rect 1796 2020 1874 2030
rect 1562 1992 1598 1994
rect 1718 1992 1754 1994
rect 1548 1986 1612 1992
rect 1548 1978 1554 1986
rect 576 1942 1554 1978
rect 576 1476 612 1942
rect 1548 1934 1554 1942
rect 1606 1934 1612 1986
rect 1548 1928 1612 1934
rect 1704 1986 1768 1992
rect 1704 1934 1710 1986
rect 1762 1934 1768 1986
rect 1796 1964 1806 2020
rect 1864 1964 1874 2020
rect 2308 1978 2348 2266
rect 2758 2260 2764 2312
rect 2816 2304 2822 2312
rect 3508 2312 3572 2318
rect 3508 2304 3514 2312
rect 2816 2268 3514 2304
rect 2816 2260 2822 2268
rect 2758 2254 2822 2260
rect 3508 2260 3514 2268
rect 3566 2260 3572 2312
rect 3638 2292 3644 2344
rect 3696 2292 3702 2344
rect 3638 2286 3702 2292
rect 3508 2254 3572 2260
rect 3522 2252 3558 2254
rect 2696 2032 2774 2042
rect 2462 1992 2498 1994
rect 2618 1992 2654 1994
rect 2448 1986 2512 1992
rect 2448 1978 2454 1986
rect 1796 1952 1874 1964
rect 2306 1940 2454 1978
rect 1704 1928 1768 1934
rect 2448 1934 2454 1940
rect 2506 1934 2512 1986
rect 2448 1928 2512 1934
rect 2604 1986 2668 1992
rect 2604 1934 2610 1986
rect 2662 1934 2668 1986
rect 2696 1976 2706 2032
rect 2764 1976 2774 2032
rect 2696 1964 2774 1976
rect 3294 2010 3372 2020
rect 3294 1954 3304 2010
rect 3362 1954 3372 2010
rect 3294 1942 3372 1954
rect 2604 1928 2668 1934
rect 1562 1926 1598 1928
rect 1718 1898 1754 1928
rect 2462 1926 2498 1928
rect 2618 1898 2654 1928
rect 884 1862 1754 1898
rect 884 1802 920 1862
rect 870 1796 934 1802
rect 870 1744 876 1796
rect 928 1744 934 1796
rect 870 1738 934 1744
rect 808 1510 886 1520
rect 562 1470 626 1476
rect 0 1458 78 1468
rect 0 1402 10 1458
rect 68 1402 78 1458
rect 562 1418 568 1470
rect 620 1418 626 1470
rect 562 1412 626 1418
rect 716 1470 780 1476
rect 716 1418 722 1470
rect 774 1418 780 1470
rect 808 1454 818 1510
rect 876 1454 886 1510
rect 808 1442 886 1454
rect 716 1412 780 1418
rect 0 1390 78 1402
rect -210 1320 62 1326
rect 576 1320 612 1412
rect -210 1284 612 1320
rect -210 1278 62 1284
rect -784 1178 -720 1184
rect -784 1126 -778 1178
rect -726 1176 -720 1178
rect -726 1152 62 1176
rect 730 1154 766 1412
rect 242 1152 766 1154
rect -726 1128 766 1152
rect -726 1126 -720 1128
rect -784 1120 -720 1126
rect 14 1116 766 1128
rect 14 1108 62 1116
rect -210 984 62 990
rect -210 948 392 984
rect -1064 934 -988 944
rect -1064 878 -1054 934
rect -998 878 -988 934
rect -1064 868 -988 878
rect -210 942 62 948
rect -778 718 -702 728
rect -778 662 -768 718
rect -712 662 -702 718
rect -778 652 -702 662
rect -1334 454 -1064 506
rect -1116 412 -1064 454
rect -1444 400 -1376 412
rect -1444 334 -1434 400
rect -1382 334 -1376 400
rect -1126 392 -1058 412
rect -1126 340 -1116 392
rect -1064 340 -1058 392
rect -1126 334 -1058 340
rect -1468 218 -1392 228
rect -1468 162 -1458 218
rect -1402 162 -1392 218
rect -1468 152 -1392 162
rect -1310 -344 -1234 -334
rect -1310 -400 -1300 -344
rect -1244 -400 -1234 -344
rect -1310 -410 -1234 -400
rect -1440 -576 -1376 -570
rect -1440 -628 -1434 -576
rect -1382 -628 -1376 -576
rect -1440 -634 -1376 -628
rect -2270 -2286 -2108 -2260
rect -2270 -2410 -2242 -2286
rect -2132 -2410 -2108 -2286
rect -2270 -2432 -2108 -2410
rect -1436 -2542 -1380 -634
rect -1340 -1368 -1276 -1362
rect -1340 -1420 -1334 -1368
rect -1282 -1420 -1276 -1368
rect -1340 -1426 -1276 -1420
rect -1334 -2448 -1282 -1426
rect -784 -1776 -720 -1770
rect -784 -1828 -778 -1776
rect -726 -1778 -720 -1776
rect -210 -1778 -162 942
rect 0 868 78 878
rect 0 812 10 868
rect 68 812 78 868
rect 0 800 78 812
rect 356 36 392 948
rect 438 114 474 1116
rect 730 996 766 1116
rect 1408 1076 1444 1862
rect 1872 1860 2654 1898
rect 1622 1778 1700 1788
rect 1622 1722 1632 1778
rect 1690 1722 1700 1778
rect 1622 1710 1700 1722
rect 1872 1416 1908 1860
rect 3652 1832 3688 2286
rect 2458 1794 3688 1832
rect 1858 1410 1922 1416
rect 1858 1358 1864 1410
rect 1916 1358 1922 1410
rect 1858 1352 1922 1358
rect 1796 1118 1874 1128
rect 1562 1090 1598 1092
rect 1718 1090 1754 1092
rect 1548 1084 1612 1090
rect 1548 1076 1554 1084
rect 1408 1040 1554 1076
rect 1548 1032 1554 1040
rect 1606 1032 1612 1084
rect 1548 1026 1612 1032
rect 1704 1084 1768 1090
rect 1704 1032 1710 1084
rect 1762 1032 1768 1084
rect 1796 1062 1806 1118
rect 1864 1062 1874 1118
rect 1796 1050 1874 1062
rect 1704 1026 1768 1032
rect 1562 1024 1598 1026
rect 1718 996 1754 1026
rect 730 960 1754 996
rect 1718 834 1754 960
rect 2458 934 2494 1794
rect 2522 1622 2600 1632
rect 2522 1566 2532 1622
rect 2590 1566 2600 1622
rect 2522 1554 2600 1566
rect 3426 1356 3504 1366
rect 3426 1300 3436 1356
rect 3494 1300 3504 1356
rect 3426 1288 3504 1300
rect 3638 1282 3702 1288
rect 2754 1254 2818 1260
rect 2754 1202 2760 1254
rect 2812 1246 2818 1254
rect 3508 1254 3572 1260
rect 3508 1246 3514 1254
rect 2812 1210 3514 1246
rect 2812 1202 2818 1210
rect 2754 1196 2818 1202
rect 3508 1202 3514 1210
rect 3566 1202 3572 1254
rect 3638 1230 3644 1282
rect 3696 1230 3702 1282
rect 3638 1224 3702 1230
rect 3508 1196 3572 1202
rect 3522 1194 3558 1196
rect 2692 968 2770 978
rect 2614 934 2650 936
rect 2444 928 2508 934
rect 2444 876 2450 928
rect 2502 876 2508 928
rect 2444 870 2508 876
rect 2600 928 2664 934
rect 2600 876 2606 928
rect 2658 876 2664 928
rect 2692 912 2702 968
rect 2760 912 2770 968
rect 2692 900 2770 912
rect 3426 948 3504 958
rect 3426 892 3436 948
rect 3494 892 3504 948
rect 3426 880 3504 892
rect 2600 870 2664 876
rect 2458 868 2494 870
rect 2614 834 2650 870
rect 634 816 712 826
rect 634 760 644 816
rect 702 760 712 816
rect 1718 798 2650 834
rect 634 748 712 760
rect 1538 550 1616 560
rect 1538 494 1548 550
rect 1606 494 1616 550
rect 3652 536 3688 1224
rect 3652 500 3902 536
rect 1538 482 1616 494
rect 1756 480 1820 486
rect 870 448 934 454
rect 870 396 876 448
rect 928 440 934 448
rect 1622 448 1686 454
rect 1622 440 1628 448
rect 928 404 1628 440
rect 928 396 934 404
rect 870 390 934 396
rect 1622 396 1628 404
rect 1680 396 1686 448
rect 1756 428 1762 480
rect 1814 472 1820 480
rect 1814 436 3902 472
rect 1814 428 1820 436
rect 1756 422 1820 428
rect 1622 390 1686 396
rect 1636 388 1672 390
rect 808 158 886 168
rect 560 122 624 128
rect 560 114 566 122
rect 438 78 566 114
rect 560 70 566 78
rect 618 70 624 122
rect 560 64 624 70
rect 716 122 780 128
rect 716 70 722 122
rect 774 70 780 122
rect 808 102 818 158
rect 876 102 886 158
rect 808 90 886 102
rect 1540 144 1618 154
rect 1540 88 1550 144
rect 1608 88 1618 144
rect 1540 76 1618 88
rect 716 64 780 70
rect 730 36 766 64
rect 356 0 766 36
rect -726 -1826 -162 -1778
rect -726 -1828 -720 -1826
rect -784 -1834 -720 -1828
rect -1064 -2020 -988 -2010
rect -1064 -2076 -1054 -2020
rect -998 -2076 -988 -2020
rect -1064 -2086 -988 -2076
rect -1068 -2168 -992 -2158
rect -1068 -2224 -1058 -2168
rect -1002 -2224 -992 -2168
rect -1068 -2234 -992 -2224
rect -778 -2356 -702 -2346
rect -778 -2412 -768 -2356
rect -712 -2412 -702 -2356
rect -778 -2422 -702 -2412
rect -1334 -2500 -1064 -2448
rect -1116 -2542 -1064 -2500
rect -1444 -2554 -1376 -2542
rect -1444 -2620 -1434 -2554
rect -1382 -2620 -1376 -2554
rect -1126 -2562 -1058 -2542
rect -1126 -2614 -1116 -2562
rect -1064 -2614 -1058 -2562
rect -1126 -2620 -1058 -2614
rect -1366 -2736 -1290 -2726
rect -1366 -2792 -1356 -2736
rect -1300 -2792 -1290 -2736
rect -1366 -2802 -1290 -2792
<< via2 >>
rect -1300 5558 -1244 5560
rect -1300 5506 -1298 5558
rect -1298 5506 -1246 5558
rect -1246 5506 -1244 5558
rect -1300 5504 -1244 5506
rect -1854 3796 -1798 3798
rect -1854 3744 -1852 3796
rect -1852 3744 -1800 3796
rect -1800 3744 -1798 3796
rect -1854 3742 -1798 3744
rect -1054 3882 -998 3884
rect -1054 3830 -1052 3882
rect -1052 3830 -1000 3882
rect -1000 3830 -998 3882
rect -1054 3828 -998 3830
rect -768 3806 -712 3808
rect -768 3754 -766 3806
rect -766 3754 -714 3806
rect -714 3754 -712 3806
rect -768 3752 -712 3754
rect -1458 3166 -1402 3168
rect -1458 3114 -1456 3166
rect -1456 3114 -1404 3166
rect -1404 3114 -1402 3166
rect -1458 3112 -1402 3114
rect -1300 2612 -1244 2614
rect -1300 2560 -1298 2612
rect -1298 2560 -1246 2612
rect -1246 2560 -1244 2612
rect -1300 2558 -1244 2560
rect 1632 2678 1690 2680
rect 1632 2626 1634 2678
rect 1634 2626 1688 2678
rect 1688 2626 1690 2678
rect 1632 2624 1690 2626
rect 2532 2678 2590 2680
rect 2532 2626 2534 2678
rect 2534 2626 2588 2678
rect 2588 2626 2590 2678
rect 2532 2624 2590 2626
rect 3436 2414 3494 2416
rect 3436 2362 3438 2414
rect 3438 2362 3492 2414
rect 3492 2362 3494 2414
rect 3436 2360 3494 2362
rect 644 2162 702 2164
rect 644 2110 646 2162
rect 646 2110 700 2162
rect 700 2110 702 2162
rect 644 2108 702 2110
rect 1806 2018 1864 2020
rect 1806 1966 1808 2018
rect 1808 1966 1862 2018
rect 1862 1966 1864 2018
rect 1806 1964 1864 1966
rect 2706 2030 2764 2032
rect 2706 1978 2708 2030
rect 2708 1978 2762 2030
rect 2762 1978 2764 2030
rect 2706 1976 2764 1978
rect 3304 2008 3362 2010
rect 3304 1956 3306 2008
rect 3306 1956 3360 2008
rect 3360 1956 3362 2008
rect 3304 1954 3362 1956
rect 10 1456 68 1458
rect 10 1404 12 1456
rect 12 1404 66 1456
rect 66 1404 68 1456
rect 10 1402 68 1404
rect 818 1508 876 1510
rect 818 1456 820 1508
rect 820 1456 874 1508
rect 874 1456 876 1508
rect 818 1454 876 1456
rect -1054 932 -998 934
rect -1054 880 -1052 932
rect -1052 880 -1000 932
rect -1000 880 -998 932
rect -1054 878 -998 880
rect -768 716 -712 718
rect -768 664 -766 716
rect -766 664 -714 716
rect -714 664 -712 716
rect -768 662 -712 664
rect -1458 216 -1402 218
rect -1458 164 -1456 216
rect -1456 164 -1404 216
rect -1404 164 -1402 216
rect -1458 162 -1402 164
rect -1300 -346 -1244 -344
rect -1300 -398 -1298 -346
rect -1298 -398 -1246 -346
rect -1246 -398 -1244 -346
rect -1300 -400 -1244 -398
rect -2242 -2410 -2132 -2286
rect 10 866 68 868
rect 10 814 12 866
rect 12 814 66 866
rect 66 814 68 866
rect 10 812 68 814
rect 1632 1776 1690 1778
rect 1632 1724 1634 1776
rect 1634 1724 1688 1776
rect 1688 1724 1690 1776
rect 1632 1722 1690 1724
rect 1806 1116 1864 1118
rect 1806 1064 1808 1116
rect 1808 1064 1862 1116
rect 1862 1064 1864 1116
rect 1806 1062 1864 1064
rect 2532 1620 2590 1622
rect 2532 1568 2534 1620
rect 2534 1568 2588 1620
rect 2588 1568 2590 1620
rect 2532 1566 2590 1568
rect 3436 1354 3494 1356
rect 3436 1302 3438 1354
rect 3438 1302 3492 1354
rect 3492 1302 3494 1354
rect 3436 1300 3494 1302
rect 2702 966 2760 968
rect 2702 914 2704 966
rect 2704 914 2758 966
rect 2758 914 2760 966
rect 2702 912 2760 914
rect 3436 946 3494 948
rect 3436 894 3438 946
rect 3438 894 3492 946
rect 3492 894 3494 946
rect 3436 892 3494 894
rect 644 814 702 816
rect 644 762 646 814
rect 646 762 700 814
rect 700 762 702 814
rect 644 760 702 762
rect 1548 548 1606 550
rect 1548 496 1550 548
rect 1550 496 1604 548
rect 1604 496 1606 548
rect 1548 494 1606 496
rect 818 156 876 158
rect 818 104 820 156
rect 820 104 874 156
rect 874 104 876 156
rect 818 102 876 104
rect 1550 142 1608 144
rect 1550 90 1552 142
rect 1552 90 1606 142
rect 1606 90 1608 142
rect 1550 88 1608 90
rect -1054 -2022 -998 -2020
rect -1054 -2074 -1052 -2022
rect -1052 -2074 -1000 -2022
rect -1000 -2074 -998 -2022
rect -1054 -2076 -998 -2074
rect -1058 -2170 -1002 -2168
rect -1058 -2222 -1056 -2170
rect -1056 -2222 -1004 -2170
rect -1004 -2222 -1002 -2170
rect -1058 -2224 -1002 -2222
rect -768 -2358 -712 -2356
rect -768 -2410 -766 -2358
rect -766 -2410 -714 -2358
rect -714 -2410 -712 -2358
rect -768 -2412 -712 -2410
rect -1356 -2738 -1300 -2736
rect -1356 -2790 -1354 -2738
rect -1354 -2790 -1302 -2738
rect -1302 -2790 -1300 -2738
rect -1356 -2792 -1300 -2790
<< metal3 >>
rect -1310 5560 -1234 5570
rect -1310 5504 -1300 5560
rect -1244 5504 -1234 5560
rect -1310 4032 -1234 5504
rect -1310 3956 -852 4032
rect -1876 3802 -1776 3820
rect -1876 3738 -1858 3802
rect -1794 3738 -1776 3802
rect -1876 3720 -1776 3738
rect -1480 3172 -1380 3190
rect -1480 3108 -1462 3172
rect -1398 3108 -1380 3172
rect -1480 3090 -1380 3108
rect -1310 2614 -1234 3956
rect -1310 2558 -1300 2614
rect -1244 2558 -1234 2614
rect -1480 222 -1380 240
rect -1480 158 -1462 222
rect -1398 158 -1380 222
rect -1480 140 -1380 158
rect -1310 -344 -1234 2558
rect -1310 -400 -1300 -344
rect -1244 -400 -1234 -344
rect -1310 -410 -1234 -400
rect -1064 3884 -988 3894
rect -1064 3828 -1054 3884
rect -998 3828 -988 3884
rect -1064 934 -988 3828
rect -928 1468 -852 3956
rect -790 3812 -690 3830
rect -790 3748 -772 3812
rect -708 3748 -690 3812
rect -790 3730 -690 3748
rect 1622 2684 1700 2690
rect 2522 2684 2600 2690
rect 1622 2680 2600 2684
rect 1622 2624 1632 2680
rect 1690 2624 2532 2680
rect 2590 2624 2600 2680
rect 1622 2620 2600 2624
rect 1622 2612 1700 2620
rect 2522 2612 2600 2620
rect 634 2168 712 2174
rect 1628 2168 1694 2612
rect 634 2164 1694 2168
rect 634 2108 644 2164
rect 702 2108 1694 2164
rect 634 2104 1694 2108
rect 634 2096 712 2104
rect -928 1462 78 1468
rect 640 1462 706 2096
rect 1628 1788 1694 2104
rect 2524 2420 2594 2612
rect 3426 2420 3504 2426
rect 2524 2416 3504 2420
rect 2524 2360 3436 2416
rect 3494 2360 3504 2416
rect 2524 2356 3504 2360
rect 1796 2020 1874 2030
rect 1796 1964 1806 2020
rect 1864 1964 1874 2020
rect 1796 1952 1874 1964
rect 1622 1778 1700 1788
rect 1622 1722 1632 1778
rect 1690 1722 1700 1778
rect 1622 1710 1700 1722
rect -928 1458 706 1462
rect -928 1402 10 1458
rect 68 1402 706 1458
rect 808 1514 886 1520
rect 1802 1514 1868 1952
rect 2524 1632 2594 2356
rect 3426 2348 3504 2356
rect 2696 2032 2774 2042
rect 2696 1976 2706 2032
rect 2764 1976 2774 2032
rect 2696 1964 2774 1976
rect 3294 2010 3372 2020
rect 2516 1622 2600 1632
rect 2516 1566 2532 1622
rect 2590 1566 2600 1622
rect 2516 1554 2600 1566
rect 808 1510 1868 1514
rect 808 1454 818 1510
rect 876 1454 1868 1510
rect 808 1450 1868 1454
rect 808 1442 886 1450
rect -928 1396 706 1402
rect -928 1390 78 1396
rect -1064 878 -1054 934
rect -998 878 -988 934
rect -1064 872 78 878
rect -1064 868 472 872
rect -1064 812 10 868
rect 68 812 472 868
rect 640 826 706 1396
rect 1802 1128 1868 1450
rect 1796 1124 1874 1128
rect 2698 1124 2768 1964
rect 3294 1954 3304 2010
rect 3362 1954 3372 2010
rect 3294 1942 3372 1954
rect 3298 1124 3368 1942
rect 3432 1366 3498 2348
rect 3428 1356 3506 1366
rect 3428 1300 3436 1356
rect 3494 1300 3506 1356
rect 3428 1288 3506 1300
rect 1796 1118 3368 1124
rect 1796 1062 1806 1118
rect 1864 1062 3368 1118
rect 1796 1058 3368 1062
rect 1796 1050 1874 1058
rect -1064 806 472 812
rect -1064 800 78 806
rect -1064 -2010 -988 800
rect -790 722 -690 740
rect -790 658 -772 722
rect -708 658 -690 722
rect -790 640 -690 658
rect 406 160 472 806
rect 634 820 712 826
rect 634 816 1610 820
rect 634 760 644 816
rect 702 760 1610 816
rect 634 756 1610 760
rect 634 748 712 756
rect 1544 560 1610 756
rect 1538 550 1616 560
rect 1538 494 1548 550
rect 1606 494 1616 550
rect 1538 482 1616 494
rect 808 160 886 168
rect 1802 160 1868 1050
rect 2698 978 2768 1058
rect 2692 968 2770 978
rect 2692 912 2702 968
rect 2760 912 2770 968
rect 2692 900 2770 912
rect 3298 958 3368 1058
rect 3298 948 3504 958
rect 3298 892 3436 948
rect 3494 892 3504 948
rect 3298 888 3504 892
rect 3426 880 3504 888
rect 406 158 1868 160
rect 406 102 818 158
rect 876 144 1868 158
rect 876 102 1550 144
rect 406 98 1550 102
rect 808 90 886 98
rect 1540 88 1550 98
rect 1608 98 1868 144
rect 1608 88 1618 98
rect 1540 76 1618 88
rect -2226 -2020 -988 -2010
rect -2226 -2076 -1054 -2020
rect -998 -2076 -988 -2020
rect -2226 -2086 -988 -2076
rect -2226 -2260 -2150 -2086
rect -1080 -2164 -980 -2146
rect -1080 -2228 -1062 -2164
rect -998 -2228 -980 -2164
rect -1080 -2246 -980 -2228
rect -2270 -2286 -2108 -2260
rect -2270 -2410 -2242 -2286
rect -2132 -2410 -2108 -2286
rect -2270 -2432 -2108 -2410
rect -790 -2352 -690 -2334
rect -790 -2416 -772 -2352
rect -708 -2416 -690 -2352
rect -790 -2434 -690 -2416
rect -1378 -2732 -1278 -2714
rect -1378 -2796 -1360 -2732
rect -1296 -2796 -1278 -2732
rect -1378 -2814 -1278 -2796
<< via3 >>
rect -1858 3798 -1794 3802
rect -1858 3742 -1854 3798
rect -1854 3742 -1798 3798
rect -1798 3742 -1794 3798
rect -1858 3738 -1794 3742
rect -1462 3168 -1398 3172
rect -1462 3112 -1458 3168
rect -1458 3112 -1402 3168
rect -1402 3112 -1398 3168
rect -1462 3108 -1398 3112
rect -1462 218 -1398 222
rect -1462 162 -1458 218
rect -1458 162 -1402 218
rect -1402 162 -1398 218
rect -1462 158 -1398 162
rect -772 3808 -708 3812
rect -772 3752 -768 3808
rect -768 3752 -712 3808
rect -712 3752 -708 3808
rect -772 3748 -708 3752
rect -772 718 -708 722
rect -772 662 -768 718
rect -768 662 -712 718
rect -712 662 -708 718
rect -772 658 -708 662
rect -1062 -2168 -998 -2164
rect -1062 -2224 -1058 -2168
rect -1058 -2224 -1002 -2168
rect -1002 -2224 -998 -2168
rect -1062 -2228 -998 -2224
rect -772 -2356 -708 -2352
rect -772 -2412 -768 -2356
rect -768 -2412 -712 -2356
rect -712 -2412 -708 -2356
rect -772 -2416 -708 -2412
rect -1360 -2736 -1296 -2732
rect -1360 -2792 -1356 -2736
rect -1356 -2792 -1300 -2736
rect -1300 -2792 -1296 -2736
rect -1360 -2796 -1296 -2792
<< metal4 >>
rect -1876 3802 -1776 3820
rect -1876 3738 -1858 3802
rect -1794 3738 -1776 3802
rect -1876 3190 -1776 3738
rect -790 3812 -690 3830
rect -790 3748 -772 3812
rect -708 3748 -690 3812
rect -1876 3172 -1380 3190
rect -1876 3108 -1462 3172
rect -1398 3108 -1380 3172
rect -1876 3090 -1380 3108
rect -1876 240 -1776 3090
rect -790 722 -690 3748
rect -790 658 -772 722
rect -708 658 -690 722
rect -1876 222 -1380 240
rect -1876 158 -1462 222
rect -1398 158 -1380 222
rect -1876 140 -1380 158
rect -1876 -2714 -1776 140
rect -790 -2146 -690 658
rect -1080 -2164 -690 -2146
rect -1080 -2228 -1062 -2164
rect -998 -2228 -690 -2164
rect -1080 -2246 -690 -2228
rect -790 -2352 -690 -2246
rect -790 -2416 -772 -2352
rect -708 -2416 -690 -2352
rect -790 -2434 -690 -2416
rect -1876 -2732 -1278 -2714
rect -1876 -2796 -1360 -2732
rect -1296 -2796 -1278 -2732
rect -1876 -2814 -1278 -2796
<< labels >>
rlabel metal1 -2268 3700 -2108 3842 1 Vref
port 4 n
rlabel metal4 -1876 3720 -1776 3820 1 Vin
port 3 n
rlabel metal4 -790 -2434 -690 -2334 5 Vbias
port 2 s
rlabel metal3 -2270 -2432 -2108 -2260 5 gnd
port 1 s
rlabel metal3 -1310 5494 -1234 5570 1 vdd
port 5 n
rlabel metal2 3862 436 3902 472 1 b1
port 6 n
rlabel metal2 3862 500 3902 536 1 b0
port 7 n
rlabel metal1 -1340 -400 -1202 -360 1 comparadorlayout_0.vdd
rlabel metal1 -1062 -2054 -990 -2010 1 comparadorlayout_0.gnd
rlabel metal1 -780 -1826 -726 -1776 1 comparadorlayout_0.out
rlabel poly -1378 -2802 -1278 -2730 5 comparadorlayout_0.Vin
rlabel poly -1220 -2802 -1120 -2730 5 comparadorlayout_0.Vref
rlabel poly -1080 -2212 -980 -2162 5 comparadorlayout_0.Vbias
rlabel metal1 -1340 2554 -1202 2594 1 comparadorlayout_1.vdd
rlabel metal1 -1062 900 -990 944 1 comparadorlayout_1.gnd
rlabel metal1 -780 1128 -726 1178 1 comparadorlayout_1.out
rlabel poly -1378 152 -1278 224 5 comparadorlayout_1.Vin
rlabel poly -1220 152 -1120 224 5 comparadorlayout_1.Vref
rlabel poly -1080 742 -980 792 5 comparadorlayout_1.Vbias
rlabel metal1 -1340 5504 -1202 5544 1 comparadorlayout_2.vdd
rlabel metal1 -1062 3850 -990 3894 1 comparadorlayout_2.gnd
rlabel metal1 -780 4078 -726 4128 1 comparadorlayout_2.out
rlabel poly -1378 3102 -1278 3174 5 comparadorlayout_2.Vin
rlabel poly -1220 3102 -1120 3174 5 comparadorlayout_2.Vref
rlabel poly -1080 3692 -980 3742 5 comparadorlayout_2.Vbias
rlabel metal2 3796 500 3832 536 1 codificador2bits_layout_0.b0
rlabel metal2 3796 436 3832 472 1 codificador2bits_layout_0.b1
rlabel metal2 20 1284 56 1320 1 codificador2bits_layout_0.c1
rlabel metal2 20 1116 56 1152 1 codificador2bits_layout_0.c2
rlabel metal2 20 948 56 984 1 codificador2bits_layout_0.c3
rlabel metal3 0 1390 78 1468 1 codificador2bits_layout_0.vdd
rlabel metal3 0 800 78 878 1 codificador2bits_layout_0.gnd
<< end >>
