magic
tech sky130A
timestamp 1702580219
<< nwell >>
rect 4115 1215 4213 1216
rect 3667 1197 3695 1202
rect 4115 1197 4145 1215
rect 3667 1185 3671 1197
rect 4115 1185 4121 1197
rect 3173 939 3201 944
rect 3173 927 3177 939
rect 3667 746 3695 751
rect 3667 734 3671 746
rect 4445 717 4468 802
rect 4445 705 4459 717
rect 4138 684 4211 689
rect 4119 668 4149 684
rect 4143 656 4149 668
<< poly >>
rect 4499 1202 4517 1203
rect 4492 1195 4524 1202
rect 4492 1178 4499 1195
rect 4517 1178 4524 1195
rect 4492 1173 4524 1178
rect 3512 1032 3544 1040
rect 3512 1015 3519 1032
rect 3537 1015 3544 1032
rect 3512 1010 3544 1015
rect 3590 1032 3622 1040
rect 3590 1015 3597 1032
rect 3615 1015 3622 1032
rect 3590 1010 3622 1015
rect 3962 1032 3994 1040
rect 3962 1015 3969 1032
rect 3987 1015 3994 1032
rect 3962 1010 3994 1015
rect 4040 1032 4072 1040
rect 4040 1015 4047 1032
rect 4065 1015 4072 1032
rect 4040 1010 4072 1015
rect 3019 774 3051 782
rect 3019 757 3026 774
rect 3044 757 3051 774
rect 3019 752 3051 757
rect 3096 774 3128 782
rect 3096 757 3103 774
rect 3121 757 3128 774
rect 3096 752 3128 757
rect 4499 673 4517 674
rect 4492 666 4524 673
rect 4492 649 4499 666
rect 4517 649 4524 666
rect 4492 644 4524 649
rect 3512 581 3544 589
rect 3512 564 3519 581
rect 3537 564 3544 581
rect 3512 559 3544 564
rect 3590 581 3622 589
rect 3590 564 3597 581
rect 3615 564 3622 581
rect 3590 559 3622 564
rect 3960 503 3992 511
rect 3960 486 3967 503
rect 3985 486 3992 503
rect 3960 481 3992 486
rect 4038 503 4070 511
rect 4038 486 4045 503
rect 4063 486 4070 503
rect 4038 481 4070 486
rect 3556 270 3574 271
rect 3549 263 3581 270
rect 3549 246 3556 263
rect 3574 246 3581 263
rect 3549 241 3581 246
<< polycont >>
rect 4499 1178 4517 1195
rect 3519 1015 3537 1032
rect 3597 1015 3615 1032
rect 3969 1015 3987 1032
rect 4047 1015 4065 1032
rect 3026 757 3044 774
rect 3103 757 3121 774
rect 4499 649 4517 666
rect 3519 564 3537 581
rect 3597 564 3615 581
rect 3967 486 3985 503
rect 4045 486 4063 503
rect 3556 246 3574 263
rect 3025 83 3043 100
rect 3103 83 3121 100
<< locali >>
rect 4499 1195 4517 1203
rect 4499 1169 4517 1178
rect 3519 1032 3537 1040
rect 3519 1006 3537 1015
rect 3597 1032 3615 1040
rect 3597 1006 3615 1015
rect 3969 1032 3987 1040
rect 3969 1006 3987 1015
rect 4047 1032 4065 1040
rect 4047 1006 4065 1015
rect 3026 774 3044 782
rect 3026 748 3044 757
rect 3103 774 3121 782
rect 3103 748 3121 757
rect 4499 666 4517 674
rect 4499 640 4517 649
rect 3519 581 3537 589
rect 3519 555 3537 564
rect 3597 581 3615 589
rect 3597 555 3615 564
rect 3967 503 3985 511
rect 3967 477 3985 486
rect 4045 503 4063 511
rect 4045 477 4063 486
rect 3556 263 3574 271
rect 3556 237 3574 246
rect 3025 100 3043 108
rect 3025 74 3043 83
rect 3103 100 3121 108
rect 3103 74 3121 83
<< viali >>
rect 4499 1178 4517 1195
rect 3519 1015 3537 1032
rect 3597 1015 3615 1032
rect 3969 1015 3987 1032
rect 4047 1015 4065 1032
rect 3026 757 3044 774
rect 3103 757 3121 774
rect 4499 649 4517 666
rect 3519 564 3537 581
rect 3597 564 3615 581
rect 3967 486 3985 503
rect 4045 486 4063 503
rect 3556 246 3574 263
rect 3025 83 3043 100
rect 3103 83 3121 100
<< metal1 >>
rect 3552 1382 3585 1385
rect 3552 1356 3555 1382
rect 3582 1356 3585 1382
rect 3552 1353 3585 1356
rect 4002 1382 4035 1385
rect 4002 1356 4005 1382
rect 4032 1356 4035 1382
rect 4002 1353 4035 1356
rect 4454 1250 4487 1253
rect 4454 1224 4457 1250
rect 4484 1224 4487 1250
rect 4454 1221 4487 1224
rect 4557 1215 4589 1218
rect 3667 1199 3699 1202
rect 3667 1173 3670 1199
rect 3696 1173 3699 1199
rect 4117 1199 4149 1202
rect 4117 1197 4120 1199
rect 4115 1175 4120 1197
rect 3667 1170 3699 1173
rect 4117 1173 4120 1175
rect 4146 1173 4149 1199
rect 4117 1170 4149 1173
rect 4492 1199 4524 1202
rect 4492 1173 4495 1199
rect 4521 1173 4524 1199
rect 4557 1189 4560 1215
rect 4586 1189 4589 1215
rect 4557 1186 4589 1189
rect 4492 1170 4524 1173
rect 3058 1124 3091 1127
rect 3058 1098 3061 1124
rect 3088 1098 3091 1124
rect 3058 1095 3091 1098
rect 4089 1058 4122 1061
rect 3639 1052 3672 1055
rect 3639 1039 3642 1052
rect 3512 1036 3544 1039
rect 3512 1010 3515 1036
rect 3541 1010 3544 1036
rect 3512 1007 3544 1010
rect 3590 1036 3622 1039
rect 3590 1010 3593 1036
rect 3619 1010 3622 1036
rect 3636 1026 3642 1039
rect 3669 1026 3672 1052
rect 3636 1023 3672 1026
rect 3962 1036 3994 1039
rect 3590 1007 3622 1010
rect 3962 1010 3965 1036
rect 3991 1010 3994 1036
rect 3962 1007 3994 1010
rect 4040 1036 4072 1039
rect 4040 1010 4043 1036
rect 4069 1010 4072 1036
rect 4089 1032 4092 1058
rect 4119 1032 4122 1058
rect 4089 1029 4122 1032
rect 4388 1049 4421 1050
rect 4388 1047 4482 1049
rect 4388 1021 4391 1047
rect 4418 1021 4482 1047
rect 4388 1019 4482 1021
rect 4388 1018 4421 1019
rect 4040 1007 4072 1010
rect 3173 941 3205 944
rect 3173 915 3176 941
rect 3202 915 3205 941
rect 3173 912 3205 915
rect 3552 931 3585 934
rect 3552 905 3555 931
rect 3582 905 3585 931
rect 3552 902 3585 905
rect 4002 853 4035 856
rect 4002 827 4005 853
rect 4032 827 4035 853
rect 4002 824 4035 827
rect 3145 797 3178 800
rect 3019 778 3051 781
rect 2741 771 2774 774
rect 2741 745 2744 771
rect 2771 745 2774 771
rect 3019 752 3022 778
rect 3048 752 3051 778
rect 3019 749 3051 752
rect 3096 778 3128 781
rect 3096 752 3099 778
rect 3125 752 3128 778
rect 3145 771 3148 797
rect 3175 771 3178 797
rect 3145 768 3178 771
rect 3096 749 3128 752
rect 2741 741 2774 745
rect 3667 748 3699 751
rect 3667 722 3670 748
rect 3696 722 3699 748
rect 3667 719 3699 722
rect 4454 720 4487 723
rect 4454 694 4457 720
rect 4484 694 4487 720
rect 4454 691 4487 694
rect 4557 684 4589 687
rect 4115 670 4147 673
rect 4115 668 4118 670
rect 4113 646 4118 668
rect 4115 644 4118 646
rect 4144 644 4147 670
rect 4115 641 4147 644
rect 4492 670 4524 673
rect 4492 644 4495 670
rect 4521 644 4524 670
rect 4557 658 4560 684
rect 4586 658 4589 684
rect 4557 655 4589 658
rect 4492 641 4524 644
rect 3639 601 3672 604
rect 3512 585 3544 588
rect 3512 559 3515 585
rect 3541 559 3544 585
rect 3512 556 3544 559
rect 3590 585 3622 588
rect 3590 559 3593 585
rect 3619 559 3622 585
rect 3639 575 3642 601
rect 3669 575 3672 601
rect 3639 572 3672 575
rect 3590 556 3622 559
rect 4087 526 4120 529
rect 3960 507 3992 510
rect 3960 481 3963 507
rect 3989 481 3992 507
rect 2741 476 2774 479
rect 3960 478 3992 481
rect 4038 507 4070 510
rect 4038 481 4041 507
rect 4067 481 4070 507
rect 4087 500 4090 526
rect 4117 500 4120 526
rect 4087 497 4120 500
rect 4454 516 4487 519
rect 4454 490 4457 516
rect 4484 490 4487 516
rect 4454 487 4487 490
rect 4038 478 4070 481
rect 2741 450 2744 476
rect 2771 450 2774 476
rect 2741 446 2774 450
rect 3058 450 3091 453
rect 3058 424 3061 450
rect 3088 424 3091 450
rect 3058 421 3091 424
rect 3510 317 3543 320
rect 3510 291 3513 317
rect 3540 291 3543 317
rect 3510 288 3543 291
rect 3616 283 3648 286
rect 3173 267 3205 270
rect 3173 265 3176 267
rect 3166 243 3176 265
rect 3173 241 3176 243
rect 3202 241 3205 267
rect 3173 238 3205 241
rect 3549 267 3581 270
rect 3549 241 3552 267
rect 3578 241 3581 267
rect 3616 257 3619 283
rect 3645 257 3648 283
rect 3616 254 3648 257
rect 3549 238 3581 241
rect 3145 121 3178 124
rect 3018 104 3050 107
rect 3018 78 3021 104
rect 3047 78 3050 104
rect 3018 75 3050 78
rect 3096 104 3128 107
rect 3096 78 3099 104
rect 3125 78 3128 104
rect 3145 95 3148 121
rect 3175 95 3178 121
rect 3145 92 3178 95
rect 3511 114 3544 117
rect 3511 88 3514 114
rect 3541 88 3544 114
rect 3511 85 3544 88
rect 3096 75 3128 78
<< via1 >>
rect 3555 1356 3582 1382
rect 4005 1356 4032 1382
rect 4457 1224 4484 1250
rect 3670 1173 3696 1199
rect 4120 1173 4146 1199
rect 4495 1195 4521 1199
rect 4495 1178 4499 1195
rect 4499 1178 4517 1195
rect 4517 1178 4521 1195
rect 4495 1173 4521 1178
rect 4560 1189 4586 1215
rect 3061 1098 3088 1124
rect 3515 1032 3541 1036
rect 3515 1015 3519 1032
rect 3519 1015 3537 1032
rect 3537 1015 3541 1032
rect 3515 1010 3541 1015
rect 3593 1032 3619 1036
rect 3593 1015 3597 1032
rect 3597 1015 3615 1032
rect 3615 1015 3619 1032
rect 3593 1010 3619 1015
rect 3642 1026 3669 1052
rect 3965 1032 3991 1036
rect 3965 1015 3969 1032
rect 3969 1015 3987 1032
rect 3987 1015 3991 1032
rect 3965 1010 3991 1015
rect 4043 1032 4069 1036
rect 4043 1015 4047 1032
rect 4047 1015 4065 1032
rect 4065 1015 4069 1032
rect 4043 1010 4069 1015
rect 4092 1032 4119 1058
rect 4391 1021 4418 1047
rect 3176 915 3202 941
rect 3555 905 3582 931
rect 4005 827 4032 853
rect 2744 745 2771 771
rect 3022 774 3048 778
rect 3022 757 3026 774
rect 3026 757 3044 774
rect 3044 757 3048 774
rect 3022 752 3048 757
rect 3099 774 3125 778
rect 3099 757 3103 774
rect 3103 757 3121 774
rect 3121 757 3125 774
rect 3099 752 3125 757
rect 3148 771 3175 797
rect 3670 722 3696 748
rect 4457 694 4484 720
rect 4118 644 4144 670
rect 4495 666 4521 670
rect 4495 649 4499 666
rect 4499 649 4517 666
rect 4517 649 4521 666
rect 4495 644 4521 649
rect 4560 658 4586 684
rect 3515 581 3541 585
rect 3515 564 3519 581
rect 3519 564 3537 581
rect 3537 564 3541 581
rect 3515 559 3541 564
rect 3593 581 3619 585
rect 3593 564 3597 581
rect 3597 564 3615 581
rect 3615 564 3619 581
rect 3593 559 3619 564
rect 3642 575 3669 601
rect 3963 503 3989 507
rect 3963 486 3967 503
rect 3967 486 3985 503
rect 3985 486 3989 503
rect 3963 481 3989 486
rect 4041 503 4067 507
rect 4041 486 4045 503
rect 4045 486 4063 503
rect 4063 486 4067 503
rect 4041 481 4067 486
rect 4090 500 4117 526
rect 4457 490 4484 516
rect 2744 450 2771 476
rect 3061 424 3088 450
rect 3513 291 3540 317
rect 3176 241 3202 267
rect 3552 263 3578 267
rect 3552 246 3556 263
rect 3556 246 3574 263
rect 3574 246 3578 263
rect 3552 241 3578 246
rect 3619 257 3645 283
rect 3021 100 3047 104
rect 3021 83 3025 100
rect 3025 83 3043 100
rect 3043 83 3047 100
rect 3021 78 3047 83
rect 3099 100 3125 104
rect 3099 83 3103 100
rect 3103 83 3121 100
rect 3121 83 3125 100
rect 3099 78 3125 83
rect 3148 95 3175 121
rect 3514 88 3541 114
<< metal2 >>
rect 3549 1383 3588 1388
rect 3549 1355 3554 1383
rect 3583 1355 3588 1383
rect 3549 1349 3588 1355
rect 3999 1383 4038 1388
rect 3999 1355 4004 1383
rect 4033 1355 4038 1383
rect 3999 1349 4038 1355
rect 4451 1251 4490 1256
rect 4451 1223 4456 1251
rect 4485 1223 4490 1251
rect 4451 1217 4490 1223
rect 4557 1215 4589 1218
rect 3667 1199 3699 1202
rect 3667 1173 3670 1199
rect 3696 1196 3699 1199
rect 4117 1199 4149 1202
rect 3696 1176 3912 1196
rect 3696 1173 3699 1176
rect 3667 1170 3699 1173
rect 3055 1125 3094 1130
rect 3055 1097 3060 1125
rect 3089 1097 3094 1125
rect 3055 1091 3094 1097
rect 3636 1053 3675 1058
rect 3519 1039 3537 1040
rect 3597 1039 3615 1040
rect 3512 1036 3544 1039
rect 3512 1032 3515 1036
rect 3026 1014 3515 1032
rect 3026 781 3044 1014
rect 3512 1010 3515 1014
rect 3541 1010 3544 1036
rect 3512 1007 3544 1010
rect 3590 1036 3622 1039
rect 3590 1010 3593 1036
rect 3619 1010 3622 1036
rect 3636 1025 3641 1053
rect 3670 1025 3675 1053
rect 3892 1032 3912 1176
rect 4117 1173 4120 1199
rect 4146 1195 4149 1199
rect 4492 1199 4524 1202
rect 4492 1195 4495 1199
rect 4146 1177 4495 1195
rect 4146 1173 4149 1177
rect 4117 1170 4149 1173
rect 4492 1173 4495 1177
rect 4521 1173 4524 1199
rect 4557 1189 4560 1215
rect 4586 1189 4589 1215
rect 4557 1186 4589 1189
rect 4492 1170 4524 1173
rect 4499 1169 4517 1170
rect 4086 1059 4125 1064
rect 3969 1039 3987 1040
rect 4047 1039 4065 1040
rect 3962 1036 3994 1039
rect 3962 1032 3965 1036
rect 3636 1019 3675 1025
rect 3891 1013 3965 1032
rect 3590 1007 3622 1010
rect 3962 1010 3965 1013
rect 3991 1010 3994 1036
rect 3962 1007 3994 1010
rect 4040 1036 4072 1039
rect 4040 1010 4043 1036
rect 4069 1010 4072 1036
rect 4086 1031 4091 1059
rect 4120 1031 4125 1059
rect 4086 1025 4125 1031
rect 4385 1048 4424 1053
rect 4385 1020 4390 1048
rect 4419 1020 4424 1048
rect 4385 1014 4424 1020
rect 4040 1007 4072 1010
rect 3519 1006 3537 1007
rect 3597 992 3615 1007
rect 3969 1006 3987 1007
rect 4047 992 4065 1007
rect 3180 974 3615 992
rect 3180 944 3198 974
rect 3173 941 3205 944
rect 3173 915 3176 941
rect 3202 915 3205 941
rect 3173 912 3205 915
rect 3142 798 3181 803
rect 3019 778 3051 781
rect 2738 772 2777 777
rect 2738 744 2743 772
rect 2772 744 2777 772
rect 3019 752 3022 778
rect 3048 752 3051 778
rect 3019 749 3051 752
rect 3096 778 3128 781
rect 3096 752 3099 778
rect 3125 752 3128 778
rect 3142 770 3147 798
rect 3176 770 3181 798
rect 3142 764 3181 770
rect 3096 749 3128 752
rect 2738 738 2777 744
rect 3026 703 3044 749
rect 2748 685 3044 703
rect 3103 620 3121 749
rect 2859 619 3121 620
rect 2748 601 3121 619
rect 2748 517 2934 535
rect 2738 477 2777 482
rect 2738 449 2743 477
rect 2772 449 2777 477
rect 2738 443 2777 449
rect 2916 61 2934 517
rect 2957 100 2975 601
rect 3103 541 3121 601
rect 3442 581 3460 974
rect 3674 973 4065 992
rect 3549 932 3588 937
rect 3549 904 3554 932
rect 3583 904 3588 932
rect 3549 898 3588 904
rect 3674 751 3692 973
rect 4564 959 4582 1186
rect 3967 940 4582 959
rect 3667 748 3699 751
rect 3667 722 3670 748
rect 3696 722 3699 748
rect 3667 719 3699 722
rect 3636 602 3675 607
rect 3519 588 3537 589
rect 3597 588 3615 589
rect 3512 585 3544 588
rect 3512 581 3515 585
rect 3442 563 3515 581
rect 3512 559 3515 563
rect 3541 559 3544 585
rect 3512 556 3544 559
rect 3590 585 3622 588
rect 3590 559 3593 585
rect 3619 559 3622 585
rect 3636 574 3641 602
rect 3670 574 3675 602
rect 3636 568 3675 574
rect 3590 556 3622 559
rect 3519 555 3537 556
rect 3597 541 3615 556
rect 3103 523 3615 541
rect 3597 460 3615 523
rect 3967 510 3985 940
rect 3999 854 4038 859
rect 3999 826 4004 854
rect 4033 826 4038 854
rect 3999 820 4038 826
rect 4451 721 4490 726
rect 4451 693 4456 721
rect 4485 693 4490 721
rect 4451 687 4490 693
rect 4557 684 4589 687
rect 4115 670 4147 673
rect 4115 644 4118 670
rect 4144 666 4147 670
rect 4492 670 4524 673
rect 4492 666 4495 670
rect 4144 648 4495 666
rect 4144 644 4147 648
rect 4115 641 4147 644
rect 4492 644 4495 648
rect 4521 644 4524 670
rect 4557 658 4560 684
rect 4586 658 4589 684
rect 4557 655 4589 658
rect 4492 641 4524 644
rect 4499 640 4517 641
rect 4084 527 4123 532
rect 4045 510 4063 511
rect 3960 507 3992 510
rect 3960 481 3963 507
rect 3989 481 3992 507
rect 3960 478 3992 481
rect 4038 507 4070 510
rect 4038 481 4041 507
rect 4067 481 4070 507
rect 4084 499 4089 527
rect 4118 499 4123 527
rect 4084 493 4123 499
rect 4451 517 4490 522
rect 4451 489 4456 517
rect 4485 489 4490 517
rect 4451 483 4490 489
rect 4038 478 4070 481
rect 3967 477 3985 478
rect 4045 460 4063 478
rect 3055 451 3094 456
rect 3055 423 3060 451
rect 3089 423 3094 451
rect 3597 442 4063 460
rect 3055 417 3094 423
rect 3507 318 3546 323
rect 3507 290 3512 318
rect 3541 290 3546 318
rect 4564 311 4582 655
rect 4564 293 4654 311
rect 3507 284 3546 290
rect 3616 283 3648 286
rect 3173 267 3205 270
rect 3173 241 3176 267
rect 3202 263 3205 267
rect 3549 267 3581 270
rect 3549 263 3552 267
rect 3202 245 3552 263
rect 3202 241 3205 245
rect 3173 238 3205 241
rect 3549 241 3552 245
rect 3578 241 3581 267
rect 3616 257 3619 283
rect 3645 279 3648 283
rect 3645 261 4654 279
rect 3645 257 3648 261
rect 3616 254 3648 257
rect 3549 238 3581 241
rect 3556 237 3574 238
rect 3142 122 3181 127
rect 3018 104 3050 107
rect 3018 100 3021 104
rect 2957 82 3021 100
rect 3018 78 3021 82
rect 3047 78 3050 104
rect 3018 75 3050 78
rect 3096 104 3128 107
rect 3096 78 3099 104
rect 3125 78 3128 104
rect 3142 94 3147 122
rect 3176 94 3181 122
rect 3142 88 3181 94
rect 3508 115 3547 120
rect 3508 87 3513 115
rect 3542 87 3547 115
rect 3508 81 3547 87
rect 3096 75 3128 78
rect 3103 61 3121 75
rect 2916 43 3121 61
<< via2 >>
rect 3554 1382 3583 1383
rect 3554 1356 3555 1382
rect 3555 1356 3582 1382
rect 3582 1356 3583 1382
rect 3554 1355 3583 1356
rect 4004 1382 4033 1383
rect 4004 1356 4005 1382
rect 4005 1356 4032 1382
rect 4032 1356 4033 1382
rect 4004 1355 4033 1356
rect 4456 1250 4485 1251
rect 4456 1224 4457 1250
rect 4457 1224 4484 1250
rect 4484 1224 4485 1250
rect 4456 1223 4485 1224
rect 3060 1124 3089 1125
rect 3060 1098 3061 1124
rect 3061 1098 3088 1124
rect 3088 1098 3089 1124
rect 3060 1097 3089 1098
rect 3641 1052 3670 1053
rect 3641 1026 3642 1052
rect 3642 1026 3669 1052
rect 3669 1026 3670 1052
rect 3641 1025 3670 1026
rect 4091 1058 4120 1059
rect 4091 1032 4092 1058
rect 4092 1032 4119 1058
rect 4119 1032 4120 1058
rect 4091 1031 4120 1032
rect 4390 1047 4419 1048
rect 4390 1021 4391 1047
rect 4391 1021 4418 1047
rect 4418 1021 4419 1047
rect 4390 1020 4419 1021
rect 2743 771 2772 772
rect 2743 745 2744 771
rect 2744 745 2771 771
rect 2771 745 2772 771
rect 2743 744 2772 745
rect 3147 797 3176 798
rect 3147 771 3148 797
rect 3148 771 3175 797
rect 3175 771 3176 797
rect 3147 770 3176 771
rect 2743 476 2772 477
rect 2743 450 2744 476
rect 2744 450 2771 476
rect 2771 450 2772 476
rect 2743 449 2772 450
rect 3554 931 3583 932
rect 3554 905 3555 931
rect 3555 905 3582 931
rect 3582 905 3583 931
rect 3554 904 3583 905
rect 3641 601 3670 602
rect 3641 575 3642 601
rect 3642 575 3669 601
rect 3669 575 3670 601
rect 3641 574 3670 575
rect 4004 853 4033 854
rect 4004 827 4005 853
rect 4005 827 4032 853
rect 4032 827 4033 853
rect 4004 826 4033 827
rect 4456 720 4485 721
rect 4456 694 4457 720
rect 4457 694 4484 720
rect 4484 694 4485 720
rect 4456 693 4485 694
rect 4089 526 4118 527
rect 4089 500 4090 526
rect 4090 500 4117 526
rect 4117 500 4118 526
rect 4089 499 4118 500
rect 4456 516 4485 517
rect 4456 490 4457 516
rect 4457 490 4484 516
rect 4484 490 4485 516
rect 4456 489 4485 490
rect 3060 450 3089 451
rect 3060 424 3061 450
rect 3061 424 3088 450
rect 3088 424 3089 450
rect 3060 423 3089 424
rect 3512 317 3541 318
rect 3512 291 3513 317
rect 3513 291 3540 317
rect 3540 291 3541 317
rect 3512 290 3541 291
rect 3147 121 3176 122
rect 3147 95 3148 121
rect 3148 95 3175 121
rect 3175 95 3176 121
rect 3147 94 3176 95
rect 3513 114 3542 115
rect 3513 88 3514 114
rect 3514 88 3541 114
rect 3541 88 3542 114
rect 3513 87 3542 88
<< metal3 >>
rect 3549 1385 3588 1388
rect 3999 1385 4038 1388
rect 3549 1383 4038 1385
rect 3549 1355 3554 1383
rect 3583 1355 4004 1383
rect 4033 1355 4038 1383
rect 3549 1353 4038 1355
rect 3549 1349 3588 1353
rect 3999 1349 4038 1353
rect 3055 1127 3094 1130
rect 3552 1127 3585 1349
rect 3055 1125 3585 1127
rect 3055 1097 3060 1125
rect 3089 1097 3585 1125
rect 3055 1095 3585 1097
rect 3055 1091 3094 1095
rect 2738 774 2777 777
rect 3058 774 3091 1091
rect 3552 937 3585 1095
rect 4000 1253 4035 1349
rect 4451 1253 4490 1256
rect 4000 1251 4490 1253
rect 4000 1223 4456 1251
rect 4485 1223 4490 1251
rect 4000 1221 4490 1223
rect 3636 1053 3675 1058
rect 3636 1025 3641 1053
rect 3670 1025 3675 1053
rect 3636 1019 3675 1025
rect 3549 932 3588 937
rect 3549 904 3554 932
rect 3583 904 3588 932
rect 3549 898 3588 904
rect 2738 772 3091 774
rect 2738 744 2743 772
rect 2772 744 3091 772
rect 3142 800 3181 803
rect 3639 800 3672 1019
rect 4000 859 4035 1221
rect 4451 1217 4490 1221
rect 4086 1059 4125 1064
rect 4086 1031 4091 1059
rect 4120 1031 4125 1059
rect 4086 1025 4125 1031
rect 4385 1048 4424 1053
rect 3996 854 4038 859
rect 3996 826 4004 854
rect 4033 826 4038 854
rect 3996 820 4038 826
rect 3142 798 3672 800
rect 3142 770 3147 798
rect 3176 770 3672 798
rect 3142 768 3672 770
rect 3142 764 3181 768
rect 2738 741 3091 744
rect 2738 738 2777 741
rect 2738 479 2777 482
rect 2738 477 2974 479
rect 2738 449 2743 477
rect 2772 449 2974 477
rect 3058 456 3091 741
rect 3639 607 3672 768
rect 3636 605 3675 607
rect 4087 605 4122 1025
rect 4385 1020 4390 1048
rect 4419 1020 4424 1048
rect 4385 1014 4424 1020
rect 4387 605 4422 1014
rect 4454 726 4487 1217
rect 4452 721 4491 726
rect 4452 693 4456 721
rect 4485 693 4491 721
rect 4452 687 4491 693
rect 3636 602 4422 605
rect 3636 574 3641 602
rect 3670 574 4422 602
rect 3636 572 4422 574
rect 3636 568 3675 572
rect 2738 446 2974 449
rect 2738 443 2777 446
rect 2941 123 2974 446
rect 3055 453 3094 456
rect 3055 451 3543 453
rect 3055 423 3060 451
rect 3089 423 3543 451
rect 3055 421 3543 423
rect 3055 417 3094 421
rect 3510 323 3543 421
rect 3507 318 3546 323
rect 3507 290 3512 318
rect 3541 290 3546 318
rect 3507 284 3546 290
rect 3142 123 3181 127
rect 3639 123 3672 568
rect 4087 532 4122 572
rect 4084 527 4123 532
rect 4084 499 4089 527
rect 4118 499 4123 527
rect 4084 493 4123 499
rect 4387 522 4422 572
rect 4387 517 4490 522
rect 4387 489 4456 517
rect 4485 489 4490 517
rect 4387 487 4490 489
rect 4451 483 4490 487
rect 2941 122 3672 123
rect 2941 94 3147 122
rect 3176 115 3672 122
rect 3176 94 3513 115
rect 2941 92 3513 94
rect 3142 88 3181 92
rect 3508 87 3513 92
rect 3542 92 3672 115
rect 3542 87 3547 92
rect 3508 81 3547 87
use nand_layout  nand_layout_0
timestamp 1702408154
transform 1 0 3341 0 1 1413
box 101 -403 422 -34
use nand_layout  nand_layout_1
timestamp 1702408154
transform 1 0 2847 0 1 481
box 101 -403 422 -34
use nand_layout  nand_layout_2
timestamp 1702408154
transform 1 0 2847 0 1 1155
box 101 -403 422 -34
use nand_layout  nand_layout_3
timestamp 1702408154
transform 1 0 3789 0 1 884
box 101 -403 422 -34
use nand_layout  nand_layout_4
timestamp 1702408154
transform 1 0 3341 0 1 962
box 101 -403 422 -34
use nand_layout  nand_layout_5
timestamp 1702408154
transform 1 0 3791 0 1 1413
box 101 -403 422 -34
use not_layout  not_layout_0
timestamp 1702580219
transform 1 0 4027 0 1 510
box 310 -20 570 333
use not_layout  not_layout_1
timestamp 1702580219
transform 1 0 3084 0 1 107
box 310 -20 570 333
use not_layout  not_layout_2
timestamp 1702580219
transform 1 0 4027 0 1 1039
box 310 -20 570 333
<< labels >>
rlabel metal2 4636 293 4654 311 1 b0
rlabel metal2 4636 261 4654 279 1 b1
rlabel metal2 2748 685 2766 703 1 c1
rlabel metal2 2748 601 2766 619 1 c2
rlabel metal2 2748 517 2766 535 1 c3
rlabel metal3 2738 738 2777 777 1 vdd
rlabel metal3 2738 443 2777 482 1 gnd
<< end >>
