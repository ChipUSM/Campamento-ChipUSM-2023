magic
tech sky130A
timestamp 1702560231
<< dnwell >>
rect -141 -2256 256 -1951
<< nwell >>
rect -176 -1091 368 -983
rect -176 -1149 300 -1091
rect -176 -1895 -92 -1149
rect 47 -1501 300 -1149
rect -176 -1979 273 -1895
rect -176 -2180 -70 -1979
rect 189 -2180 273 -1979
rect -176 -2264 273 -2180
<< pwell >>
rect -70 -2180 189 -1979
<< mvnmos >>
rect 74 -1827 124 -1727
rect 218 -1827 268 -1785
rect -5 -2121 45 -2071
rect 74 -2121 124 -2071
<< mvpmos >>
rect -114 -1066 -64 -1016
rect -35 -1066 15 -1016
rect 109 -1468 159 -1018
rect 188 -1468 238 -1018
<< mvndiff >>
rect 45 -1733 74 -1727
rect 45 -1821 51 -1733
rect 68 -1821 74 -1733
rect 45 -1827 74 -1821
rect 124 -1733 153 -1727
rect 124 -1821 130 -1733
rect 147 -1821 153 -1733
rect 124 -1827 153 -1821
rect 189 -1791 218 -1785
rect 189 -1821 195 -1791
rect 212 -1821 218 -1791
rect 189 -1827 218 -1821
rect 268 -1791 297 -1785
rect 268 -1821 274 -1791
rect 291 -1821 297 -1791
rect 268 -1827 297 -1821
rect -34 -2077 -5 -2071
rect -34 -2115 -28 -2077
rect -11 -2115 -5 -2077
rect -34 -2121 -5 -2115
rect 45 -2077 74 -2071
rect 45 -2115 51 -2077
rect 68 -2115 74 -2077
rect 45 -2121 74 -2115
rect 124 -2077 153 -2071
rect 124 -2115 130 -2077
rect 147 -2115 153 -2077
rect 124 -2121 153 -2115
<< mvpdiff >>
rect -143 -1022 -114 -1016
rect -143 -1060 -137 -1022
rect -120 -1060 -114 -1022
rect -143 -1066 -114 -1060
rect -64 -1022 -35 -1016
rect -64 -1060 -58 -1022
rect -41 -1060 -35 -1022
rect -64 -1066 -35 -1060
rect 15 -1022 44 -1016
rect 15 -1060 21 -1022
rect 38 -1060 44 -1022
rect 15 -1066 44 -1060
rect 80 -1024 109 -1018
rect 80 -1462 86 -1024
rect 103 -1462 109 -1024
rect 80 -1468 109 -1462
rect 159 -1024 188 -1018
rect 159 -1462 165 -1024
rect 182 -1462 188 -1024
rect 159 -1468 188 -1462
rect 238 -1024 267 -1018
rect 238 -1462 244 -1024
rect 261 -1462 267 -1024
rect 238 -1468 267 -1462
<< mvndiffc >>
rect 51 -1821 68 -1733
rect 130 -1821 147 -1733
rect 195 -1821 212 -1791
rect 274 -1821 291 -1791
rect -28 -2115 -11 -2077
rect 51 -2115 68 -2077
rect 130 -2115 147 -2077
<< mvpdiffc >>
rect -137 -1060 -120 -1022
rect -58 -1060 -41 -1022
rect 21 -1060 38 -1022
rect 86 -1462 103 -1024
rect 165 -1462 182 -1024
rect 244 -1462 261 -1024
<< mvpsubdiff >>
rect 118 -1666 159 -1661
rect 118 -1685 130 -1666
rect 147 -1685 159 -1666
rect 118 -1690 159 -1685
rect 39 -1996 80 -1992
rect 39 -2031 51 -1996
rect 68 -2031 80 -1996
rect 39 -2034 80 -2031
<< mvnsubdiff >>
rect 294 -1028 335 -1016
rect 294 -1046 306 -1028
rect 323 -1046 335 -1028
rect 294 -1058 335 -1046
<< mvpsubdiffcont >>
rect 130 -1685 147 -1666
rect 51 -2031 68 -1996
<< mvnsubdiffcont >>
rect 306 -1046 323 -1028
<< poly >>
rect -114 -1016 -64 -1003
rect -35 -1016 15 -1003
rect 109 -1018 159 -1005
rect 188 -1018 238 -1005
rect -114 -1079 -64 -1066
rect -35 -1079 15 -1066
rect -143 -1091 15 -1079
rect -143 -1110 -137 -1091
rect -120 -1110 -30 -1091
rect -143 -1111 -30 -1110
rect -10 -1111 15 -1091
rect -143 -1123 15 -1111
rect 109 -1479 159 -1468
rect 188 -1479 238 -1468
rect 80 -1493 238 -1479
rect 80 -1510 97 -1493
rect 120 -1510 238 -1493
rect 80 -1523 238 -1510
rect 74 -1727 124 -1714
rect 218 -1785 268 -1772
rect 74 -1840 124 -1827
rect 218 -1840 268 -1827
rect 74 -1881 268 -1840
rect 144 -1906 194 -1881
rect -5 -2071 45 -2058
rect 74 -2071 124 -2058
rect -5 -2201 45 -2121
rect 74 -2201 124 -2121
<< polycont >>
rect -137 -1110 -120 -1091
rect -30 -1111 -10 -1091
rect 97 -1510 120 -1493
<< locali >>
rect -137 -1022 -120 -1014
rect -137 -1091 -120 -1060
rect -58 -1022 -41 -1014
rect -58 -1068 -41 -1060
rect 21 -1022 38 -1014
rect 21 -1068 38 -1060
rect 86 -1024 103 -1016
rect -137 -1118 -120 -1110
rect -30 -1091 -10 -1083
rect -30 -1119 -10 -1111
rect 86 -1470 103 -1462
rect 165 -1024 182 -1016
rect 165 -1470 182 -1462
rect 244 -1024 261 -1016
rect 306 -1028 323 -1018
rect 261 -1046 306 -1028
rect 306 -1056 323 -1046
rect 244 -1470 261 -1462
rect 20 -1487 40 -1481
rect 20 -1513 40 -1507
rect 89 -1510 97 -1493
rect 120 -1510 128 -1493
rect 130 -1666 147 -1654
rect 51 -1733 68 -1725
rect 51 -1829 68 -1821
rect 130 -1733 147 -1685
rect 130 -1829 147 -1821
rect 195 -1791 212 -1783
rect 195 -1829 212 -1821
rect 274 -1791 291 -1783
rect 274 -1829 291 -1821
rect 51 -1996 68 -1988
rect -28 -2077 -11 -2069
rect -28 -2123 -11 -2115
rect 51 -2077 68 -2031
rect 51 -2123 68 -2115
rect 130 -2077 147 -2069
rect 130 -2123 147 -2115
<< viali >>
rect -137 -1060 -120 -1022
rect -58 -1060 -41 -1022
rect 21 -1060 38 -1022
rect -30 -1111 -10 -1091
rect 86 -1462 103 -1024
rect 165 -1462 182 -1024
rect 244 -1462 261 -1024
rect 20 -1507 40 -1487
rect 97 -1510 120 -1493
rect 51 -1821 68 -1733
rect 130 -1821 147 -1733
rect 195 -1821 212 -1791
rect 274 -1821 291 -1791
rect -28 -2115 -11 -2077
rect 51 -2115 68 -2077
rect 130 -2115 147 -2077
<< metal1 >>
rect -61 -1000 264 -980
rect -140 -1022 -117 -1016
rect -140 -1060 -137 -1022
rect -120 -1060 -117 -1022
rect -140 -1066 -117 -1060
rect -61 -1022 -38 -1000
rect -61 -1060 -58 -1022
rect -41 -1060 -38 -1022
rect -61 -1066 -38 -1060
rect 18 -1022 41 -1016
rect 18 -1060 21 -1022
rect 38 -1060 41 -1022
rect -36 -1088 -4 -1085
rect -36 -1114 -33 -1088
rect -7 -1114 -4 -1088
rect -36 -1117 -4 -1114
rect 18 -1481 41 -1060
rect 83 -1024 106 -1000
rect 83 -1462 86 -1024
rect 103 -1462 106 -1024
rect 83 -1468 106 -1462
rect 162 -1024 185 -1018
rect 162 -1462 165 -1024
rect 182 -1462 185 -1024
rect 14 -1484 46 -1481
rect 14 -1510 17 -1484
rect 43 -1490 46 -1484
rect 43 -1493 126 -1490
rect 43 -1510 97 -1493
rect 120 -1510 126 -1493
rect 14 -1513 126 -1510
rect 162 -1688 185 -1462
rect 241 -1024 264 -1000
rect 241 -1462 244 -1024
rect 261 -1462 264 -1024
rect 241 -1468 264 -1462
rect 162 -1713 321 -1688
rect 48 -1733 71 -1727
rect 48 -1821 51 -1733
rect 68 -1821 71 -1733
rect -38 -2077 -4 -2071
rect -38 -2110 -33 -2077
rect -7 -2110 -4 -2077
rect 48 -2077 71 -1821
rect 127 -1733 150 -1727
rect 127 -1821 130 -1733
rect 147 -1805 150 -1733
rect 192 -1791 215 -1785
rect 192 -1805 195 -1791
rect 147 -1821 195 -1805
rect 212 -1821 215 -1791
rect 127 -1827 215 -1821
rect 271 -1791 294 -1713
rect 271 -1821 274 -1791
rect 291 -1821 294 -1791
rect 271 -1827 294 -1821
rect -31 -2115 -28 -2110
rect -11 -2115 -8 -2110
rect -31 -2121 -8 -2115
rect 48 -2115 51 -2077
rect 68 -2115 71 -2077
rect 121 -2077 155 -2071
rect 121 -2081 130 -2077
rect 147 -2081 155 -2077
rect 121 -2107 126 -2081
rect 152 -2107 155 -2081
rect 121 -2110 130 -2107
rect 48 -2121 71 -2115
rect 127 -2115 130 -2110
rect 147 -2110 155 -2107
rect 147 -2115 150 -2110
rect 127 -2121 150 -2115
<< via1 >>
rect -33 -1091 -7 -1088
rect -33 -1111 -30 -1091
rect -30 -1111 -10 -1091
rect -10 -1111 -7 -1091
rect -33 -1114 -7 -1111
rect 17 -1487 43 -1484
rect 17 -1507 20 -1487
rect 20 -1507 40 -1487
rect 40 -1507 43 -1487
rect 17 -1510 43 -1507
rect -33 -2110 -28 -2077
rect -28 -2110 -11 -2077
rect -11 -2110 -7 -2077
rect 126 -2107 130 -2081
rect 130 -2107 147 -2081
rect 147 -2107 152 -2081
<< metal2 >>
rect -36 -1088 -4 -1085
rect -36 -1114 -33 -1088
rect -7 -1114 -4 -1088
rect -36 -1117 -4 -1114
rect -34 -2071 -6 -1117
rect 14 -1484 46 -1481
rect 14 -1510 17 -1484
rect 43 -1510 46 -1484
rect 14 -1513 46 -1510
rect 17 -2024 43 -1513
rect 17 -2050 152 -2024
rect 126 -2071 152 -2050
rect -38 -2077 -4 -2071
rect -38 -2110 -33 -2077
rect -7 -2110 -4 -2077
rect 121 -2081 155 -2071
rect 121 -2107 126 -2081
rect 152 -2107 155 -2081
rect 121 -2110 155 -2107
<< labels >>
rlabel metal1 14 -1000 83 -980 1 vdd
port 1 n
rlabel metal1 153 -1827 189 -1805 1 gnd
port 2 n
rlabel metal1 294 -1713 321 -1688 1 out
port 3 n
rlabel poly -5 -2201 45 -2165 5 Vin
port 4 s
rlabel poly 74 -2201 124 -2165 5 Vref
port 5 s
rlabel poly 144 -1906 194 -1881 5 Vbias
port 6 s
<< end >>
