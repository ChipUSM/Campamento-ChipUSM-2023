magic
tech sky130A
magscale 1 2
timestamp 1702410929
<< poly >>
rect -35 777 35 793
rect -35 743 -19 777
rect 19 743 35 777
rect -35 363 35 743
rect -35 -743 35 -363
rect -35 -777 -19 -743
rect 19 -777 35 -743
rect -35 -793 35 -777
<< polycont >>
rect -19 743 19 777
rect -19 -777 19 -743
<< npolyres >>
rect -35 -363 35 363
<< locali >>
rect -35 743 -19 777
rect 19 743 35 777
rect -35 -777 -19 -743
rect 19 -777 35 -743
<< viali >>
rect -19 743 19 777
rect -19 380 19 743
rect -19 -743 19 -380
rect -19 -777 19 -743
<< metal1 >>
rect -25 777 25 789
rect -25 380 -19 777
rect 19 380 25 777
rect -25 368 25 380
rect -25 -380 25 -368
rect -25 -777 -19 -380
rect 19 -777 25 -380
rect -25 -789 25 -777
<< properties >>
string gencell sky130_fd_pr__res_generic_po
string library sky130
string parameters w 0.35 l 3.631 m 1 nx 1 wmin 0.330 lmin 1.650 rho 48.2 val 500.04 dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 0 guard 0 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 hv_guard 0 n_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
