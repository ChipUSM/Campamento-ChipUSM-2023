magic
tech sky130A
magscale 1 2
timestamp 1702434633
<< xpolycontact >>
rect -285 124 285 556
rect -285 -556 285 -124
<< xpolyres >>
rect -285 -124 285 124
<< viali >>
rect -269 141 269 538
rect -269 -538 269 -141
<< metal1 >>
rect -281 538 281 544
rect -281 141 -269 538
rect 269 141 281 538
rect -281 135 281 141
rect -281 -141 281 -135
rect -281 -538 -269 -141
rect 269 -538 281 -141
rect -281 -544 281 -538
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_2p85
string library sky130
string parameters w 2.85 l 1.237 m 1 nx 1 wmin 2.850 lmin 0.50 rho 2000 val 1.0k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 2.850 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
