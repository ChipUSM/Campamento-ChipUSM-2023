magic
tech sky130A
magscale 1 2
timestamp 1702434633
<< xpolycontact >>
rect -285 52 285 484
rect -285 -484 285 -52
<< xpolyres >>
rect -285 -52 285 52
<< viali >>
rect -269 69 269 466
rect -269 -466 269 -69
<< metal1 >>
rect -281 466 281 472
rect -281 69 -269 466
rect 269 69 281 466
rect -281 63 281 69
rect -281 -69 281 -63
rect -281 -466 -269 -69
rect 269 -466 281 -69
rect -281 -472 281 -466
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_2p85
string library sky130
string parameters w 2.85 l 0.524 m 1 nx 1 wmin 2.850 lmin 0.50 rho 2000 val 499.789 dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 2.850 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
